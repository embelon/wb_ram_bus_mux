VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_ram_bus_mux
  CLASS BLOCK ;
  FOREIGN wb_ram_bus_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 400.000 ;
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 12.875 10.640 14.475 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.195 10.640 30.795 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.515 10.640 47.115 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.035 10.640 22.635 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.355 10.640 38.955 389.200 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END wb_rst_i
  PIN wbs_hr_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 219.000 60.000 219.600 ;
    END
  END wbs_hr_ack_i
  PIN wbs_hr_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 8.200 60.000 8.800 ;
    END
  END wbs_hr_cyc_o
  PIN wbs_hr_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 224.440 60.000 225.040 ;
    END
  END wbs_hr_dat_i[0]
  PIN wbs_hr_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 280.200 60.000 280.800 ;
    END
  END wbs_hr_dat_i[10]
  PIN wbs_hr_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 285.640 60.000 286.240 ;
    END
  END wbs_hr_dat_i[11]
  PIN wbs_hr_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 291.080 60.000 291.680 ;
    END
  END wbs_hr_dat_i[12]
  PIN wbs_hr_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 296.520 60.000 297.120 ;
    END
  END wbs_hr_dat_i[13]
  PIN wbs_hr_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 302.640 60.000 303.240 ;
    END
  END wbs_hr_dat_i[14]
  PIN wbs_hr_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 308.080 60.000 308.680 ;
    END
  END wbs_hr_dat_i[15]
  PIN wbs_hr_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 313.520 60.000 314.120 ;
    END
  END wbs_hr_dat_i[16]
  PIN wbs_hr_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 318.960 60.000 319.560 ;
    END
  END wbs_hr_dat_i[17]
  PIN wbs_hr_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 324.400 60.000 325.000 ;
    END
  END wbs_hr_dat_i[18]
  PIN wbs_hr_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 329.840 60.000 330.440 ;
    END
  END wbs_hr_dat_i[19]
  PIN wbs_hr_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 229.880 60.000 230.480 ;
    END
  END wbs_hr_dat_i[1]
  PIN wbs_hr_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 335.960 60.000 336.560 ;
    END
  END wbs_hr_dat_i[20]
  PIN wbs_hr_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 341.400 60.000 342.000 ;
    END
  END wbs_hr_dat_i[21]
  PIN wbs_hr_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 346.840 60.000 347.440 ;
    END
  END wbs_hr_dat_i[22]
  PIN wbs_hr_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 352.280 60.000 352.880 ;
    END
  END wbs_hr_dat_i[23]
  PIN wbs_hr_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 357.720 60.000 358.320 ;
    END
  END wbs_hr_dat_i[24]
  PIN wbs_hr_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 363.160 60.000 363.760 ;
    END
  END wbs_hr_dat_i[25]
  PIN wbs_hr_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 369.280 60.000 369.880 ;
    END
  END wbs_hr_dat_i[26]
  PIN wbs_hr_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 374.720 60.000 375.320 ;
    END
  END wbs_hr_dat_i[27]
  PIN wbs_hr_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 380.160 60.000 380.760 ;
    END
  END wbs_hr_dat_i[28]
  PIN wbs_hr_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 385.600 60.000 386.200 ;
    END
  END wbs_hr_dat_i[29]
  PIN wbs_hr_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 236.000 60.000 236.600 ;
    END
  END wbs_hr_dat_i[2]
  PIN wbs_hr_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 391.040 60.000 391.640 ;
    END
  END wbs_hr_dat_i[30]
  PIN wbs_hr_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 396.480 60.000 397.080 ;
    END
  END wbs_hr_dat_i[31]
  PIN wbs_hr_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 241.440 60.000 242.040 ;
    END
  END wbs_hr_dat_i[3]
  PIN wbs_hr_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 246.880 60.000 247.480 ;
    END
  END wbs_hr_dat_i[4]
  PIN wbs_hr_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 252.320 60.000 252.920 ;
    END
  END wbs_hr_dat_i[5]
  PIN wbs_hr_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 257.760 60.000 258.360 ;
    END
  END wbs_hr_dat_i[6]
  PIN wbs_hr_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 263.200 60.000 263.800 ;
    END
  END wbs_hr_dat_i[7]
  PIN wbs_hr_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 269.320 60.000 269.920 ;
    END
  END wbs_hr_dat_i[8]
  PIN wbs_hr_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 274.760 60.000 275.360 ;
    END
  END wbs_hr_dat_i[9]
  PIN wbs_hr_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 41.520 60.000 42.120 ;
    END
  END wbs_hr_dat_o[0]
  PIN wbs_hr_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 96.600 60.000 97.200 ;
    END
  END wbs_hr_dat_o[10]
  PIN wbs_hr_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 102.720 60.000 103.320 ;
    END
  END wbs_hr_dat_o[11]
  PIN wbs_hr_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 108.160 60.000 108.760 ;
    END
  END wbs_hr_dat_o[12]
  PIN wbs_hr_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 113.600 60.000 114.200 ;
    END
  END wbs_hr_dat_o[13]
  PIN wbs_hr_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 119.040 60.000 119.640 ;
    END
  END wbs_hr_dat_o[14]
  PIN wbs_hr_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 124.480 60.000 125.080 ;
    END
  END wbs_hr_dat_o[15]
  PIN wbs_hr_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 129.920 60.000 130.520 ;
    END
  END wbs_hr_dat_o[16]
  PIN wbs_hr_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 136.040 60.000 136.640 ;
    END
  END wbs_hr_dat_o[17]
  PIN wbs_hr_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 141.480 60.000 142.080 ;
    END
  END wbs_hr_dat_o[18]
  PIN wbs_hr_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 146.920 60.000 147.520 ;
    END
  END wbs_hr_dat_o[19]
  PIN wbs_hr_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 46.960 60.000 47.560 ;
    END
  END wbs_hr_dat_o[1]
  PIN wbs_hr_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 152.360 60.000 152.960 ;
    END
  END wbs_hr_dat_o[20]
  PIN wbs_hr_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 157.800 60.000 158.400 ;
    END
  END wbs_hr_dat_o[21]
  PIN wbs_hr_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 163.240 60.000 163.840 ;
    END
  END wbs_hr_dat_o[22]
  PIN wbs_hr_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 169.360 60.000 169.960 ;
    END
  END wbs_hr_dat_o[23]
  PIN wbs_hr_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 174.800 60.000 175.400 ;
    END
  END wbs_hr_dat_o[24]
  PIN wbs_hr_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 180.240 60.000 180.840 ;
    END
  END wbs_hr_dat_o[25]
  PIN wbs_hr_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 185.680 60.000 186.280 ;
    END
  END wbs_hr_dat_o[26]
  PIN wbs_hr_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 191.120 60.000 191.720 ;
    END
  END wbs_hr_dat_o[27]
  PIN wbs_hr_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 196.560 60.000 197.160 ;
    END
  END wbs_hr_dat_o[28]
  PIN wbs_hr_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 202.680 60.000 203.280 ;
    END
  END wbs_hr_dat_o[29]
  PIN wbs_hr_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 52.400 60.000 53.000 ;
    END
  END wbs_hr_dat_o[2]
  PIN wbs_hr_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 208.120 60.000 208.720 ;
    END
  END wbs_hr_dat_o[30]
  PIN wbs_hr_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 213.560 60.000 214.160 ;
    END
  END wbs_hr_dat_o[31]
  PIN wbs_hr_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 57.840 60.000 58.440 ;
    END
  END wbs_hr_dat_o[3]
  PIN wbs_hr_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 63.280 60.000 63.880 ;
    END
  END wbs_hr_dat_o[4]
  PIN wbs_hr_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 69.400 60.000 70.000 ;
    END
  END wbs_hr_dat_o[5]
  PIN wbs_hr_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 74.840 60.000 75.440 ;
    END
  END wbs_hr_dat_o[6]
  PIN wbs_hr_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 80.280 60.000 80.880 ;
    END
  END wbs_hr_dat_o[7]
  PIN wbs_hr_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 85.720 60.000 86.320 ;
    END
  END wbs_hr_dat_o[8]
  PIN wbs_hr_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 91.160 60.000 91.760 ;
    END
  END wbs_hr_dat_o[9]
  PIN wbs_hr_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 19.080 60.000 19.680 ;
    END
  END wbs_hr_sel_o[0]
  PIN wbs_hr_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 24.520 60.000 25.120 ;
    END
  END wbs_hr_sel_o[1]
  PIN wbs_hr_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 29.960 60.000 30.560 ;
    END
  END wbs_hr_sel_o[2]
  PIN wbs_hr_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 36.080 60.000 36.680 ;
    END
  END wbs_hr_sel_o[3]
  PIN wbs_hr_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 2.760 60.000 3.360 ;
    END
  END wbs_hr_stb_o
  PIN wbs_hr_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 13.640 60.000 14.240 ;
    END
  END wbs_hr_we_o
  PIN wbs_or_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END wbs_or_ack_i
  PIN wbs_or_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END wbs_or_cyc_o
  PIN wbs_or_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END wbs_or_dat_i[0]
  PIN wbs_or_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END wbs_or_dat_i[10]
  PIN wbs_or_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END wbs_or_dat_i[11]
  PIN wbs_or_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END wbs_or_dat_i[12]
  PIN wbs_or_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END wbs_or_dat_i[13]
  PIN wbs_or_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END wbs_or_dat_i[14]
  PIN wbs_or_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END wbs_or_dat_i[15]
  PIN wbs_or_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END wbs_or_dat_i[16]
  PIN wbs_or_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END wbs_or_dat_i[17]
  PIN wbs_or_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END wbs_or_dat_i[18]
  PIN wbs_or_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END wbs_or_dat_i[19]
  PIN wbs_or_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END wbs_or_dat_i[1]
  PIN wbs_or_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END wbs_or_dat_i[20]
  PIN wbs_or_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END wbs_or_dat_i[21]
  PIN wbs_or_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END wbs_or_dat_i[22]
  PIN wbs_or_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END wbs_or_dat_i[23]
  PIN wbs_or_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END wbs_or_dat_i[24]
  PIN wbs_or_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END wbs_or_dat_i[25]
  PIN wbs_or_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END wbs_or_dat_i[26]
  PIN wbs_or_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END wbs_or_dat_i[27]
  PIN wbs_or_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END wbs_or_dat_i[28]
  PIN wbs_or_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END wbs_or_dat_i[29]
  PIN wbs_or_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END wbs_or_dat_i[2]
  PIN wbs_or_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END wbs_or_dat_i[30]
  PIN wbs_or_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END wbs_or_dat_i[31]
  PIN wbs_or_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END wbs_or_dat_i[3]
  PIN wbs_or_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END wbs_or_dat_i[4]
  PIN wbs_or_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END wbs_or_dat_i[5]
  PIN wbs_or_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END wbs_or_dat_i[6]
  PIN wbs_or_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END wbs_or_dat_i[7]
  PIN wbs_or_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END wbs_or_dat_i[8]
  PIN wbs_or_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END wbs_or_dat_i[9]
  PIN wbs_or_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END wbs_or_dat_o[0]
  PIN wbs_or_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END wbs_or_dat_o[10]
  PIN wbs_or_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END wbs_or_dat_o[11]
  PIN wbs_or_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END wbs_or_dat_o[12]
  PIN wbs_or_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END wbs_or_dat_o[13]
  PIN wbs_or_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END wbs_or_dat_o[14]
  PIN wbs_or_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END wbs_or_dat_o[15]
  PIN wbs_or_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END wbs_or_dat_o[16]
  PIN wbs_or_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END wbs_or_dat_o[17]
  PIN wbs_or_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END wbs_or_dat_o[18]
  PIN wbs_or_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END wbs_or_dat_o[19]
  PIN wbs_or_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END wbs_or_dat_o[1]
  PIN wbs_or_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END wbs_or_dat_o[20]
  PIN wbs_or_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END wbs_or_dat_o[21]
  PIN wbs_or_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END wbs_or_dat_o[22]
  PIN wbs_or_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END wbs_or_dat_o[23]
  PIN wbs_or_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END wbs_or_dat_o[24]
  PIN wbs_or_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END wbs_or_dat_o[25]
  PIN wbs_or_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END wbs_or_dat_o[26]
  PIN wbs_or_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END wbs_or_dat_o[27]
  PIN wbs_or_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END wbs_or_dat_o[28]
  PIN wbs_or_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END wbs_or_dat_o[29]
  PIN wbs_or_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END wbs_or_dat_o[2]
  PIN wbs_or_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END wbs_or_dat_o[30]
  PIN wbs_or_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END wbs_or_dat_o[31]
  PIN wbs_or_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END wbs_or_dat_o[3]
  PIN wbs_or_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END wbs_or_dat_o[4]
  PIN wbs_or_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END wbs_or_dat_o[5]
  PIN wbs_or_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END wbs_or_dat_o[6]
  PIN wbs_or_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END wbs_or_dat_o[7]
  PIN wbs_or_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END wbs_or_dat_o[8]
  PIN wbs_or_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END wbs_or_dat_o[9]
  PIN wbs_or_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END wbs_or_sel_o[0]
  PIN wbs_or_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END wbs_or_sel_o[1]
  PIN wbs_or_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END wbs_or_sel_o[2]
  PIN wbs_or_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END wbs_or_sel_o[3]
  PIN wbs_or_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END wbs_or_stb_o
  PIN wbs_or_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END wbs_or_we_o
  PIN wbs_ufp_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END wbs_ufp_ack_o
  PIN wbs_ufp_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END wbs_ufp_adr_i[0]
  PIN wbs_ufp_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END wbs_ufp_adr_i[10]
  PIN wbs_ufp_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END wbs_ufp_adr_i[11]
  PIN wbs_ufp_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wbs_ufp_adr_i[12]
  PIN wbs_ufp_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END wbs_ufp_adr_i[13]
  PIN wbs_ufp_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END wbs_ufp_adr_i[14]
  PIN wbs_ufp_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wbs_ufp_adr_i[15]
  PIN wbs_ufp_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END wbs_ufp_adr_i[16]
  PIN wbs_ufp_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END wbs_ufp_adr_i[17]
  PIN wbs_ufp_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END wbs_ufp_adr_i[18]
  PIN wbs_ufp_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END wbs_ufp_adr_i[19]
  PIN wbs_ufp_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END wbs_ufp_adr_i[1]
  PIN wbs_ufp_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END wbs_ufp_adr_i[20]
  PIN wbs_ufp_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END wbs_ufp_adr_i[21]
  PIN wbs_ufp_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END wbs_ufp_adr_i[22]
  PIN wbs_ufp_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END wbs_ufp_adr_i[23]
  PIN wbs_ufp_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wbs_ufp_adr_i[24]
  PIN wbs_ufp_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END wbs_ufp_adr_i[25]
  PIN wbs_ufp_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END wbs_ufp_adr_i[26]
  PIN wbs_ufp_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END wbs_ufp_adr_i[27]
  PIN wbs_ufp_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END wbs_ufp_adr_i[28]
  PIN wbs_ufp_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END wbs_ufp_adr_i[29]
  PIN wbs_ufp_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END wbs_ufp_adr_i[2]
  PIN wbs_ufp_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END wbs_ufp_adr_i[30]
  PIN wbs_ufp_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END wbs_ufp_adr_i[31]
  PIN wbs_ufp_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wbs_ufp_adr_i[3]
  PIN wbs_ufp_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END wbs_ufp_adr_i[4]
  PIN wbs_ufp_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END wbs_ufp_adr_i[5]
  PIN wbs_ufp_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END wbs_ufp_adr_i[6]
  PIN wbs_ufp_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END wbs_ufp_adr_i[7]
  PIN wbs_ufp_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END wbs_ufp_adr_i[8]
  PIN wbs_ufp_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END wbs_ufp_adr_i[9]
  PIN wbs_ufp_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END wbs_ufp_cyc_i
  PIN wbs_ufp_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END wbs_ufp_dat_i[0]
  PIN wbs_ufp_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END wbs_ufp_dat_i[10]
  PIN wbs_ufp_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END wbs_ufp_dat_i[11]
  PIN wbs_ufp_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END wbs_ufp_dat_i[12]
  PIN wbs_ufp_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END wbs_ufp_dat_i[13]
  PIN wbs_ufp_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END wbs_ufp_dat_i[14]
  PIN wbs_ufp_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END wbs_ufp_dat_i[15]
  PIN wbs_ufp_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END wbs_ufp_dat_i[16]
  PIN wbs_ufp_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END wbs_ufp_dat_i[17]
  PIN wbs_ufp_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END wbs_ufp_dat_i[18]
  PIN wbs_ufp_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END wbs_ufp_dat_i[19]
  PIN wbs_ufp_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END wbs_ufp_dat_i[1]
  PIN wbs_ufp_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wbs_ufp_dat_i[20]
  PIN wbs_ufp_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END wbs_ufp_dat_i[21]
  PIN wbs_ufp_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END wbs_ufp_dat_i[22]
  PIN wbs_ufp_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END wbs_ufp_dat_i[23]
  PIN wbs_ufp_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END wbs_ufp_dat_i[24]
  PIN wbs_ufp_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END wbs_ufp_dat_i[25]
  PIN wbs_ufp_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END wbs_ufp_dat_i[26]
  PIN wbs_ufp_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END wbs_ufp_dat_i[27]
  PIN wbs_ufp_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END wbs_ufp_dat_i[28]
  PIN wbs_ufp_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END wbs_ufp_dat_i[29]
  PIN wbs_ufp_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END wbs_ufp_dat_i[2]
  PIN wbs_ufp_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END wbs_ufp_dat_i[30]
  PIN wbs_ufp_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END wbs_ufp_dat_i[31]
  PIN wbs_ufp_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END wbs_ufp_dat_i[3]
  PIN wbs_ufp_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END wbs_ufp_dat_i[4]
  PIN wbs_ufp_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END wbs_ufp_dat_i[5]
  PIN wbs_ufp_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END wbs_ufp_dat_i[6]
  PIN wbs_ufp_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END wbs_ufp_dat_i[7]
  PIN wbs_ufp_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END wbs_ufp_dat_i[8]
  PIN wbs_ufp_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END wbs_ufp_dat_i[9]
  PIN wbs_ufp_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END wbs_ufp_dat_o[0]
  PIN wbs_ufp_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END wbs_ufp_dat_o[10]
  PIN wbs_ufp_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END wbs_ufp_dat_o[11]
  PIN wbs_ufp_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END wbs_ufp_dat_o[12]
  PIN wbs_ufp_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END wbs_ufp_dat_o[13]
  PIN wbs_ufp_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END wbs_ufp_dat_o[14]
  PIN wbs_ufp_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END wbs_ufp_dat_o[15]
  PIN wbs_ufp_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END wbs_ufp_dat_o[16]
  PIN wbs_ufp_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END wbs_ufp_dat_o[17]
  PIN wbs_ufp_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END wbs_ufp_dat_o[18]
  PIN wbs_ufp_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END wbs_ufp_dat_o[19]
  PIN wbs_ufp_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END wbs_ufp_dat_o[1]
  PIN wbs_ufp_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END wbs_ufp_dat_o[20]
  PIN wbs_ufp_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END wbs_ufp_dat_o[21]
  PIN wbs_ufp_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END wbs_ufp_dat_o[22]
  PIN wbs_ufp_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END wbs_ufp_dat_o[23]
  PIN wbs_ufp_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END wbs_ufp_dat_o[24]
  PIN wbs_ufp_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END wbs_ufp_dat_o[25]
  PIN wbs_ufp_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END wbs_ufp_dat_o[26]
  PIN wbs_ufp_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END wbs_ufp_dat_o[27]
  PIN wbs_ufp_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END wbs_ufp_dat_o[28]
  PIN wbs_ufp_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END wbs_ufp_dat_o[29]
  PIN wbs_ufp_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END wbs_ufp_dat_o[2]
  PIN wbs_ufp_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END wbs_ufp_dat_o[30]
  PIN wbs_ufp_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END wbs_ufp_dat_o[31]
  PIN wbs_ufp_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END wbs_ufp_dat_o[3]
  PIN wbs_ufp_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END wbs_ufp_dat_o[4]
  PIN wbs_ufp_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END wbs_ufp_dat_o[5]
  PIN wbs_ufp_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END wbs_ufp_dat_o[6]
  PIN wbs_ufp_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END wbs_ufp_dat_o[7]
  PIN wbs_ufp_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END wbs_ufp_dat_o[8]
  PIN wbs_ufp_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END wbs_ufp_dat_o[9]
  PIN wbs_ufp_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END wbs_ufp_sel_i[0]
  PIN wbs_ufp_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END wbs_ufp_sel_i[1]
  PIN wbs_ufp_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END wbs_ufp_sel_i[2]
  PIN wbs_ufp_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END wbs_ufp_sel_i[3]
  PIN wbs_ufp_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END wbs_ufp_stb_i
  PIN wbs_ufp_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END wbs_ufp_we_i
  OBS
      LAYER li1 ;
        RECT 1.065 3.145 55.515 391.255 ;
      LAYER met1 ;
        RECT 0.070 3.100 55.575 391.300 ;
      LAYER met2 ;
        RECT 0.100 2.875 55.110 398.325 ;
      LAYER met3 ;
        RECT 4.400 397.480 56.000 398.305 ;
        RECT 4.400 397.440 55.600 397.480 ;
        RECT 4.000 396.800 55.600 397.440 ;
        RECT 4.400 396.080 55.600 396.800 ;
        RECT 4.400 395.400 56.000 396.080 ;
        RECT 4.000 394.760 56.000 395.400 ;
        RECT 4.400 393.360 56.000 394.760 ;
        RECT 4.000 392.040 56.000 393.360 ;
        RECT 4.400 390.640 55.600 392.040 ;
        RECT 4.000 390.000 56.000 390.640 ;
        RECT 4.400 388.600 56.000 390.000 ;
        RECT 4.000 387.960 56.000 388.600 ;
        RECT 4.400 386.600 56.000 387.960 ;
        RECT 4.400 386.560 55.600 386.600 ;
        RECT 4.000 385.240 55.600 386.560 ;
        RECT 4.400 385.200 55.600 385.240 ;
        RECT 4.400 383.840 56.000 385.200 ;
        RECT 4.000 383.200 56.000 383.840 ;
        RECT 4.400 381.800 56.000 383.200 ;
        RECT 4.000 381.160 56.000 381.800 ;
        RECT 4.400 379.760 55.600 381.160 ;
        RECT 4.000 378.440 56.000 379.760 ;
        RECT 4.400 377.040 56.000 378.440 ;
        RECT 4.000 376.400 56.000 377.040 ;
        RECT 4.400 375.720 56.000 376.400 ;
        RECT 4.400 375.000 55.600 375.720 ;
        RECT 4.000 374.360 55.600 375.000 ;
        RECT 4.400 374.320 55.600 374.360 ;
        RECT 4.400 372.960 56.000 374.320 ;
        RECT 4.000 372.320 56.000 372.960 ;
        RECT 4.400 370.920 56.000 372.320 ;
        RECT 4.000 370.280 56.000 370.920 ;
        RECT 4.000 369.600 55.600 370.280 ;
        RECT 4.400 368.880 55.600 369.600 ;
        RECT 4.400 368.200 56.000 368.880 ;
        RECT 4.000 367.560 56.000 368.200 ;
        RECT 4.400 366.160 56.000 367.560 ;
        RECT 4.000 365.520 56.000 366.160 ;
        RECT 4.400 364.160 56.000 365.520 ;
        RECT 4.400 364.120 55.600 364.160 ;
        RECT 4.000 362.800 55.600 364.120 ;
        RECT 4.400 362.760 55.600 362.800 ;
        RECT 4.400 361.400 56.000 362.760 ;
        RECT 4.000 360.760 56.000 361.400 ;
        RECT 4.400 359.360 56.000 360.760 ;
        RECT 4.000 358.720 56.000 359.360 ;
        RECT 4.400 357.320 55.600 358.720 ;
        RECT 4.000 356.000 56.000 357.320 ;
        RECT 4.400 354.600 56.000 356.000 ;
        RECT 4.000 353.960 56.000 354.600 ;
        RECT 4.400 353.280 56.000 353.960 ;
        RECT 4.400 352.560 55.600 353.280 ;
        RECT 4.000 351.920 55.600 352.560 ;
        RECT 4.400 351.880 55.600 351.920 ;
        RECT 4.400 350.520 56.000 351.880 ;
        RECT 4.000 349.880 56.000 350.520 ;
        RECT 4.400 348.480 56.000 349.880 ;
        RECT 4.000 347.840 56.000 348.480 ;
        RECT 4.000 347.160 55.600 347.840 ;
        RECT 4.400 346.440 55.600 347.160 ;
        RECT 4.400 345.760 56.000 346.440 ;
        RECT 4.000 345.120 56.000 345.760 ;
        RECT 4.400 343.720 56.000 345.120 ;
        RECT 4.000 343.080 56.000 343.720 ;
        RECT 4.400 342.400 56.000 343.080 ;
        RECT 4.400 341.680 55.600 342.400 ;
        RECT 4.000 341.000 55.600 341.680 ;
        RECT 4.000 340.360 56.000 341.000 ;
        RECT 4.400 338.960 56.000 340.360 ;
        RECT 4.000 338.320 56.000 338.960 ;
        RECT 4.400 336.960 56.000 338.320 ;
        RECT 4.400 336.920 55.600 336.960 ;
        RECT 4.000 336.280 55.600 336.920 ;
        RECT 4.400 335.560 55.600 336.280 ;
        RECT 4.400 334.880 56.000 335.560 ;
        RECT 4.000 333.560 56.000 334.880 ;
        RECT 4.400 332.160 56.000 333.560 ;
        RECT 4.000 331.520 56.000 332.160 ;
        RECT 4.400 330.840 56.000 331.520 ;
        RECT 4.400 330.120 55.600 330.840 ;
        RECT 4.000 329.480 55.600 330.120 ;
        RECT 4.400 329.440 55.600 329.480 ;
        RECT 4.400 328.080 56.000 329.440 ;
        RECT 4.000 326.760 56.000 328.080 ;
        RECT 4.400 325.400 56.000 326.760 ;
        RECT 4.400 325.360 55.600 325.400 ;
        RECT 4.000 324.720 55.600 325.360 ;
        RECT 4.400 324.000 55.600 324.720 ;
        RECT 4.400 323.320 56.000 324.000 ;
        RECT 4.000 322.680 56.000 323.320 ;
        RECT 4.400 321.280 56.000 322.680 ;
        RECT 4.000 320.640 56.000 321.280 ;
        RECT 4.400 319.960 56.000 320.640 ;
        RECT 4.400 319.240 55.600 319.960 ;
        RECT 4.000 318.560 55.600 319.240 ;
        RECT 4.000 317.920 56.000 318.560 ;
        RECT 4.400 316.520 56.000 317.920 ;
        RECT 4.000 315.880 56.000 316.520 ;
        RECT 4.400 314.520 56.000 315.880 ;
        RECT 4.400 314.480 55.600 314.520 ;
        RECT 4.000 313.840 55.600 314.480 ;
        RECT 4.400 313.120 55.600 313.840 ;
        RECT 4.400 312.440 56.000 313.120 ;
        RECT 4.000 311.120 56.000 312.440 ;
        RECT 4.400 309.720 56.000 311.120 ;
        RECT 4.000 309.080 56.000 309.720 ;
        RECT 4.400 307.680 55.600 309.080 ;
        RECT 4.000 307.040 56.000 307.680 ;
        RECT 4.400 305.640 56.000 307.040 ;
        RECT 4.000 304.320 56.000 305.640 ;
        RECT 4.400 303.640 56.000 304.320 ;
        RECT 4.400 302.920 55.600 303.640 ;
        RECT 4.000 302.280 55.600 302.920 ;
        RECT 4.400 302.240 55.600 302.280 ;
        RECT 4.400 300.880 56.000 302.240 ;
        RECT 4.000 300.240 56.000 300.880 ;
        RECT 4.400 298.840 56.000 300.240 ;
        RECT 4.000 298.200 56.000 298.840 ;
        RECT 4.400 297.520 56.000 298.200 ;
        RECT 4.400 296.800 55.600 297.520 ;
        RECT 4.000 296.120 55.600 296.800 ;
        RECT 4.000 295.480 56.000 296.120 ;
        RECT 4.400 294.080 56.000 295.480 ;
        RECT 4.000 293.440 56.000 294.080 ;
        RECT 4.400 292.080 56.000 293.440 ;
        RECT 4.400 292.040 55.600 292.080 ;
        RECT 4.000 291.400 55.600 292.040 ;
        RECT 4.400 290.680 55.600 291.400 ;
        RECT 4.400 290.000 56.000 290.680 ;
        RECT 4.000 288.680 56.000 290.000 ;
        RECT 4.400 287.280 56.000 288.680 ;
        RECT 4.000 286.640 56.000 287.280 ;
        RECT 4.400 285.240 55.600 286.640 ;
        RECT 4.000 284.600 56.000 285.240 ;
        RECT 4.400 283.200 56.000 284.600 ;
        RECT 4.000 281.880 56.000 283.200 ;
        RECT 4.400 281.200 56.000 281.880 ;
        RECT 4.400 280.480 55.600 281.200 ;
        RECT 4.000 279.840 55.600 280.480 ;
        RECT 4.400 279.800 55.600 279.840 ;
        RECT 4.400 278.440 56.000 279.800 ;
        RECT 4.000 277.800 56.000 278.440 ;
        RECT 4.400 276.400 56.000 277.800 ;
        RECT 4.000 275.760 56.000 276.400 ;
        RECT 4.400 274.360 55.600 275.760 ;
        RECT 4.000 273.040 56.000 274.360 ;
        RECT 4.400 271.640 56.000 273.040 ;
        RECT 4.000 271.000 56.000 271.640 ;
        RECT 4.400 270.320 56.000 271.000 ;
        RECT 4.400 269.600 55.600 270.320 ;
        RECT 4.000 268.960 55.600 269.600 ;
        RECT 4.400 268.920 55.600 268.960 ;
        RECT 4.400 267.560 56.000 268.920 ;
        RECT 4.000 266.240 56.000 267.560 ;
        RECT 4.400 264.840 56.000 266.240 ;
        RECT 4.000 264.200 56.000 264.840 ;
        RECT 4.400 262.800 55.600 264.200 ;
        RECT 4.000 262.160 56.000 262.800 ;
        RECT 4.400 260.760 56.000 262.160 ;
        RECT 4.000 259.440 56.000 260.760 ;
        RECT 4.400 258.760 56.000 259.440 ;
        RECT 4.400 258.040 55.600 258.760 ;
        RECT 4.000 257.400 55.600 258.040 ;
        RECT 4.400 257.360 55.600 257.400 ;
        RECT 4.400 256.000 56.000 257.360 ;
        RECT 4.000 255.360 56.000 256.000 ;
        RECT 4.400 253.960 56.000 255.360 ;
        RECT 4.000 253.320 56.000 253.960 ;
        RECT 4.000 252.640 55.600 253.320 ;
        RECT 4.400 251.920 55.600 252.640 ;
        RECT 4.400 251.240 56.000 251.920 ;
        RECT 4.000 250.600 56.000 251.240 ;
        RECT 4.400 249.200 56.000 250.600 ;
        RECT 4.000 248.560 56.000 249.200 ;
        RECT 4.400 247.880 56.000 248.560 ;
        RECT 4.400 247.160 55.600 247.880 ;
        RECT 4.000 246.520 55.600 247.160 ;
        RECT 4.400 246.480 55.600 246.520 ;
        RECT 4.400 245.120 56.000 246.480 ;
        RECT 4.000 243.800 56.000 245.120 ;
        RECT 4.400 242.440 56.000 243.800 ;
        RECT 4.400 242.400 55.600 242.440 ;
        RECT 4.000 241.760 55.600 242.400 ;
        RECT 4.400 241.040 55.600 241.760 ;
        RECT 4.400 240.360 56.000 241.040 ;
        RECT 4.000 239.720 56.000 240.360 ;
        RECT 4.400 238.320 56.000 239.720 ;
        RECT 4.000 237.000 56.000 238.320 ;
        RECT 4.400 235.600 55.600 237.000 ;
        RECT 4.000 234.960 56.000 235.600 ;
        RECT 4.400 233.560 56.000 234.960 ;
        RECT 4.000 232.920 56.000 233.560 ;
        RECT 4.400 231.520 56.000 232.920 ;
        RECT 4.000 230.880 56.000 231.520 ;
        RECT 4.000 230.200 55.600 230.880 ;
        RECT 4.400 229.480 55.600 230.200 ;
        RECT 4.400 228.800 56.000 229.480 ;
        RECT 4.000 228.160 56.000 228.800 ;
        RECT 4.400 226.760 56.000 228.160 ;
        RECT 4.000 226.120 56.000 226.760 ;
        RECT 4.400 225.440 56.000 226.120 ;
        RECT 4.400 224.720 55.600 225.440 ;
        RECT 4.000 224.080 55.600 224.720 ;
        RECT 4.400 224.040 55.600 224.080 ;
        RECT 4.400 222.680 56.000 224.040 ;
        RECT 4.000 221.360 56.000 222.680 ;
        RECT 4.400 220.000 56.000 221.360 ;
        RECT 4.400 219.960 55.600 220.000 ;
        RECT 4.000 219.320 55.600 219.960 ;
        RECT 4.400 218.600 55.600 219.320 ;
        RECT 4.400 217.920 56.000 218.600 ;
        RECT 4.000 217.280 56.000 217.920 ;
        RECT 4.400 215.880 56.000 217.280 ;
        RECT 4.000 214.560 56.000 215.880 ;
        RECT 4.400 213.160 55.600 214.560 ;
        RECT 4.000 212.520 56.000 213.160 ;
        RECT 4.400 211.120 56.000 212.520 ;
        RECT 4.000 210.480 56.000 211.120 ;
        RECT 4.400 209.120 56.000 210.480 ;
        RECT 4.400 209.080 55.600 209.120 ;
        RECT 4.000 207.760 55.600 209.080 ;
        RECT 4.400 207.720 55.600 207.760 ;
        RECT 4.400 206.360 56.000 207.720 ;
        RECT 4.000 205.720 56.000 206.360 ;
        RECT 4.400 204.320 56.000 205.720 ;
        RECT 4.000 203.680 56.000 204.320 ;
        RECT 4.400 202.280 55.600 203.680 ;
        RECT 4.000 201.640 56.000 202.280 ;
        RECT 4.400 200.240 56.000 201.640 ;
        RECT 4.000 198.920 56.000 200.240 ;
        RECT 4.400 197.560 56.000 198.920 ;
        RECT 4.400 197.520 55.600 197.560 ;
        RECT 4.000 196.880 55.600 197.520 ;
        RECT 4.400 196.160 55.600 196.880 ;
        RECT 4.400 195.480 56.000 196.160 ;
        RECT 4.000 194.840 56.000 195.480 ;
        RECT 4.400 193.440 56.000 194.840 ;
        RECT 4.000 192.120 56.000 193.440 ;
        RECT 4.400 190.720 55.600 192.120 ;
        RECT 4.000 190.080 56.000 190.720 ;
        RECT 4.400 188.680 56.000 190.080 ;
        RECT 4.000 188.040 56.000 188.680 ;
        RECT 4.400 186.680 56.000 188.040 ;
        RECT 4.400 186.640 55.600 186.680 ;
        RECT 4.000 185.320 55.600 186.640 ;
        RECT 4.400 185.280 55.600 185.320 ;
        RECT 4.400 183.920 56.000 185.280 ;
        RECT 4.000 183.280 56.000 183.920 ;
        RECT 4.400 181.880 56.000 183.280 ;
        RECT 4.000 181.240 56.000 181.880 ;
        RECT 4.400 179.840 55.600 181.240 ;
        RECT 4.000 178.520 56.000 179.840 ;
        RECT 4.400 177.120 56.000 178.520 ;
        RECT 4.000 176.480 56.000 177.120 ;
        RECT 4.400 175.800 56.000 176.480 ;
        RECT 4.400 175.080 55.600 175.800 ;
        RECT 4.000 174.440 55.600 175.080 ;
        RECT 4.400 174.400 55.600 174.440 ;
        RECT 4.400 173.040 56.000 174.400 ;
        RECT 4.000 172.400 56.000 173.040 ;
        RECT 4.400 171.000 56.000 172.400 ;
        RECT 4.000 170.360 56.000 171.000 ;
        RECT 4.000 169.680 55.600 170.360 ;
        RECT 4.400 168.960 55.600 169.680 ;
        RECT 4.400 168.280 56.000 168.960 ;
        RECT 4.000 167.640 56.000 168.280 ;
        RECT 4.400 166.240 56.000 167.640 ;
        RECT 4.000 165.600 56.000 166.240 ;
        RECT 4.400 164.240 56.000 165.600 ;
        RECT 4.400 164.200 55.600 164.240 ;
        RECT 4.000 162.880 55.600 164.200 ;
        RECT 4.400 162.840 55.600 162.880 ;
        RECT 4.400 161.480 56.000 162.840 ;
        RECT 4.000 160.840 56.000 161.480 ;
        RECT 4.400 159.440 56.000 160.840 ;
        RECT 4.000 158.800 56.000 159.440 ;
        RECT 4.400 157.400 55.600 158.800 ;
        RECT 4.000 156.080 56.000 157.400 ;
        RECT 4.400 154.680 56.000 156.080 ;
        RECT 4.000 154.040 56.000 154.680 ;
        RECT 4.400 153.360 56.000 154.040 ;
        RECT 4.400 152.640 55.600 153.360 ;
        RECT 4.000 152.000 55.600 152.640 ;
        RECT 4.400 151.960 55.600 152.000 ;
        RECT 4.400 150.600 56.000 151.960 ;
        RECT 4.000 149.960 56.000 150.600 ;
        RECT 4.400 148.560 56.000 149.960 ;
        RECT 4.000 147.920 56.000 148.560 ;
        RECT 4.000 147.240 55.600 147.920 ;
        RECT 4.400 146.520 55.600 147.240 ;
        RECT 4.400 145.840 56.000 146.520 ;
        RECT 4.000 145.200 56.000 145.840 ;
        RECT 4.400 143.800 56.000 145.200 ;
        RECT 4.000 143.160 56.000 143.800 ;
        RECT 4.400 142.480 56.000 143.160 ;
        RECT 4.400 141.760 55.600 142.480 ;
        RECT 4.000 141.080 55.600 141.760 ;
        RECT 4.000 140.440 56.000 141.080 ;
        RECT 4.400 139.040 56.000 140.440 ;
        RECT 4.000 138.400 56.000 139.040 ;
        RECT 4.400 137.040 56.000 138.400 ;
        RECT 4.400 137.000 55.600 137.040 ;
        RECT 4.000 136.360 55.600 137.000 ;
        RECT 4.400 135.640 55.600 136.360 ;
        RECT 4.400 134.960 56.000 135.640 ;
        RECT 4.000 133.640 56.000 134.960 ;
        RECT 4.400 132.240 56.000 133.640 ;
        RECT 4.000 131.600 56.000 132.240 ;
        RECT 4.400 130.920 56.000 131.600 ;
        RECT 4.400 130.200 55.600 130.920 ;
        RECT 4.000 129.560 55.600 130.200 ;
        RECT 4.400 129.520 55.600 129.560 ;
        RECT 4.400 128.160 56.000 129.520 ;
        RECT 4.000 126.840 56.000 128.160 ;
        RECT 4.400 125.480 56.000 126.840 ;
        RECT 4.400 125.440 55.600 125.480 ;
        RECT 4.000 124.800 55.600 125.440 ;
        RECT 4.400 124.080 55.600 124.800 ;
        RECT 4.400 123.400 56.000 124.080 ;
        RECT 4.000 122.760 56.000 123.400 ;
        RECT 4.400 121.360 56.000 122.760 ;
        RECT 4.000 120.720 56.000 121.360 ;
        RECT 4.400 120.040 56.000 120.720 ;
        RECT 4.400 119.320 55.600 120.040 ;
        RECT 4.000 118.640 55.600 119.320 ;
        RECT 4.000 118.000 56.000 118.640 ;
        RECT 4.400 116.600 56.000 118.000 ;
        RECT 4.000 115.960 56.000 116.600 ;
        RECT 4.400 114.600 56.000 115.960 ;
        RECT 4.400 114.560 55.600 114.600 ;
        RECT 4.000 113.920 55.600 114.560 ;
        RECT 4.400 113.200 55.600 113.920 ;
        RECT 4.400 112.520 56.000 113.200 ;
        RECT 4.000 111.200 56.000 112.520 ;
        RECT 4.400 109.800 56.000 111.200 ;
        RECT 4.000 109.160 56.000 109.800 ;
        RECT 4.400 107.760 55.600 109.160 ;
        RECT 4.000 107.120 56.000 107.760 ;
        RECT 4.400 105.720 56.000 107.120 ;
        RECT 4.000 104.400 56.000 105.720 ;
        RECT 4.400 103.720 56.000 104.400 ;
        RECT 4.400 103.000 55.600 103.720 ;
        RECT 4.000 102.360 55.600 103.000 ;
        RECT 4.400 102.320 55.600 102.360 ;
        RECT 4.400 100.960 56.000 102.320 ;
        RECT 4.000 100.320 56.000 100.960 ;
        RECT 4.400 98.920 56.000 100.320 ;
        RECT 4.000 98.280 56.000 98.920 ;
        RECT 4.400 97.600 56.000 98.280 ;
        RECT 4.400 96.880 55.600 97.600 ;
        RECT 4.000 96.200 55.600 96.880 ;
        RECT 4.000 95.560 56.000 96.200 ;
        RECT 4.400 94.160 56.000 95.560 ;
        RECT 4.000 93.520 56.000 94.160 ;
        RECT 4.400 92.160 56.000 93.520 ;
        RECT 4.400 92.120 55.600 92.160 ;
        RECT 4.000 91.480 55.600 92.120 ;
        RECT 4.400 90.760 55.600 91.480 ;
        RECT 4.400 90.080 56.000 90.760 ;
        RECT 4.000 88.760 56.000 90.080 ;
        RECT 4.400 87.360 56.000 88.760 ;
        RECT 4.000 86.720 56.000 87.360 ;
        RECT 4.400 85.320 55.600 86.720 ;
        RECT 4.000 84.680 56.000 85.320 ;
        RECT 4.400 83.280 56.000 84.680 ;
        RECT 4.000 81.960 56.000 83.280 ;
        RECT 4.400 81.280 56.000 81.960 ;
        RECT 4.400 80.560 55.600 81.280 ;
        RECT 4.000 79.920 55.600 80.560 ;
        RECT 4.400 79.880 55.600 79.920 ;
        RECT 4.400 78.520 56.000 79.880 ;
        RECT 4.000 77.880 56.000 78.520 ;
        RECT 4.400 76.480 56.000 77.880 ;
        RECT 4.000 75.840 56.000 76.480 ;
        RECT 4.400 74.440 55.600 75.840 ;
        RECT 4.000 73.120 56.000 74.440 ;
        RECT 4.400 71.720 56.000 73.120 ;
        RECT 4.000 71.080 56.000 71.720 ;
        RECT 4.400 70.400 56.000 71.080 ;
        RECT 4.400 69.680 55.600 70.400 ;
        RECT 4.000 69.040 55.600 69.680 ;
        RECT 4.400 69.000 55.600 69.040 ;
        RECT 4.400 67.640 56.000 69.000 ;
        RECT 4.000 66.320 56.000 67.640 ;
        RECT 4.400 64.920 56.000 66.320 ;
        RECT 4.000 64.280 56.000 64.920 ;
        RECT 4.400 62.880 55.600 64.280 ;
        RECT 4.000 62.240 56.000 62.880 ;
        RECT 4.400 60.840 56.000 62.240 ;
        RECT 4.000 59.520 56.000 60.840 ;
        RECT 4.400 58.840 56.000 59.520 ;
        RECT 4.400 58.120 55.600 58.840 ;
        RECT 4.000 57.480 55.600 58.120 ;
        RECT 4.400 57.440 55.600 57.480 ;
        RECT 4.400 56.080 56.000 57.440 ;
        RECT 4.000 55.440 56.000 56.080 ;
        RECT 4.400 54.040 56.000 55.440 ;
        RECT 4.000 53.400 56.000 54.040 ;
        RECT 4.000 52.720 55.600 53.400 ;
        RECT 4.400 52.000 55.600 52.720 ;
        RECT 4.400 51.320 56.000 52.000 ;
        RECT 4.000 50.680 56.000 51.320 ;
        RECT 4.400 49.280 56.000 50.680 ;
        RECT 4.000 48.640 56.000 49.280 ;
        RECT 4.400 47.960 56.000 48.640 ;
        RECT 4.400 47.240 55.600 47.960 ;
        RECT 4.000 46.600 55.600 47.240 ;
        RECT 4.400 46.560 55.600 46.600 ;
        RECT 4.400 45.200 56.000 46.560 ;
        RECT 4.000 43.880 56.000 45.200 ;
        RECT 4.400 42.520 56.000 43.880 ;
        RECT 4.400 42.480 55.600 42.520 ;
        RECT 4.000 41.840 55.600 42.480 ;
        RECT 4.400 41.120 55.600 41.840 ;
        RECT 4.400 40.440 56.000 41.120 ;
        RECT 4.000 39.800 56.000 40.440 ;
        RECT 4.400 38.400 56.000 39.800 ;
        RECT 4.000 37.080 56.000 38.400 ;
        RECT 4.400 35.680 55.600 37.080 ;
        RECT 4.000 35.040 56.000 35.680 ;
        RECT 4.400 33.640 56.000 35.040 ;
        RECT 4.000 33.000 56.000 33.640 ;
        RECT 4.400 31.600 56.000 33.000 ;
        RECT 4.000 30.960 56.000 31.600 ;
        RECT 4.000 30.280 55.600 30.960 ;
        RECT 4.400 29.560 55.600 30.280 ;
        RECT 4.400 28.880 56.000 29.560 ;
        RECT 4.000 28.240 56.000 28.880 ;
        RECT 4.400 26.840 56.000 28.240 ;
        RECT 4.000 26.200 56.000 26.840 ;
        RECT 4.400 25.520 56.000 26.200 ;
        RECT 4.400 24.800 55.600 25.520 ;
        RECT 4.000 24.160 55.600 24.800 ;
        RECT 4.400 24.120 55.600 24.160 ;
        RECT 4.400 22.760 56.000 24.120 ;
        RECT 4.000 21.440 56.000 22.760 ;
        RECT 4.400 20.080 56.000 21.440 ;
        RECT 4.400 20.040 55.600 20.080 ;
        RECT 4.000 19.400 55.600 20.040 ;
        RECT 4.400 18.680 55.600 19.400 ;
        RECT 4.400 18.000 56.000 18.680 ;
        RECT 4.000 17.360 56.000 18.000 ;
        RECT 4.400 15.960 56.000 17.360 ;
        RECT 4.000 14.640 56.000 15.960 ;
        RECT 4.400 13.240 55.600 14.640 ;
        RECT 4.000 12.600 56.000 13.240 ;
        RECT 4.400 11.200 56.000 12.600 ;
        RECT 4.000 10.560 56.000 11.200 ;
        RECT 4.400 9.200 56.000 10.560 ;
        RECT 4.400 9.160 55.600 9.200 ;
        RECT 4.000 7.840 55.600 9.160 ;
        RECT 4.400 7.800 55.600 7.840 ;
        RECT 4.400 6.440 56.000 7.800 ;
        RECT 4.000 5.800 56.000 6.440 ;
        RECT 4.400 4.400 56.000 5.800 ;
        RECT 4.000 3.760 56.000 4.400 ;
        RECT 4.400 2.895 55.600 3.760 ;
      LAYER met4 ;
        RECT 5.815 10.640 12.475 389.200 ;
        RECT 14.875 10.640 20.635 389.200 ;
        RECT 23.035 10.640 28.795 389.200 ;
        RECT 31.195 10.640 33.745 389.200 ;
  END
END wb_ram_bus_mux
END LIBRARY

