magic
tech sky130A
magscale 1 2
timestamp 1636582060
<< locali >>
rect 10977 77027 11011 78217
rect 765 49351 799 53533
rect 857 51051 891 52309
rect 949 52139 983 60809
rect 949 50847 983 51765
rect 857 50813 983 50847
rect 213 46087 247 46733
rect 857 42279 891 50813
rect 949 44795 983 48297
rect 10977 44523 11011 48501
rect 11069 44795 11103 47413
rect 857 36091 891 42109
rect 949 36839 983 43061
rect 10977 18751 11011 21369
rect 10977 14399 11011 17561
rect 11069 12835 11103 17289
rect 3617 5559 3651 5797
rect 10977 3043 11011 5593
rect 10977 663 11011 2805
rect 11069 2431 11103 5865
<< viali >>
rect 10977 78217 11011 78251
rect 1409 77469 1443 77503
rect 2053 77469 2087 77503
rect 2881 77469 2915 77503
rect 3985 77469 4019 77503
rect 9505 77469 9539 77503
rect 10149 77469 10183 77503
rect 1593 77333 1627 77367
rect 2237 77333 2271 77367
rect 2697 77333 2731 77367
rect 3801 77333 3835 77367
rect 9321 77333 9355 77367
rect 9965 77333 9999 77367
rect 1409 76993 1443 77027
rect 2053 76993 2087 77027
rect 2881 76993 2915 77027
rect 10149 76993 10183 77027
rect 10977 76993 11011 77027
rect 1593 76789 1627 76823
rect 2237 76789 2271 76823
rect 2697 76789 2731 76823
rect 9965 76789 9999 76823
rect 1409 76381 1443 76415
rect 2237 76381 2271 76415
rect 2697 76381 2731 76415
rect 10149 76381 10183 76415
rect 1593 76245 1627 76279
rect 2053 76245 2087 76279
rect 2881 76245 2915 76279
rect 9965 76245 9999 76279
rect 1593 76041 1627 76075
rect 2053 76041 2087 76075
rect 1409 75905 1443 75939
rect 2237 75905 2271 75939
rect 1777 75429 1811 75463
rect 1956 75293 1990 75327
rect 2053 75293 2087 75327
rect 2329 75293 2363 75327
rect 2789 75293 2823 75327
rect 10149 75293 10183 75327
rect 2145 75225 2179 75259
rect 2973 75157 3007 75191
rect 9965 75157 9999 75191
rect 3157 74885 3191 74919
rect 3249 74885 3283 74919
rect 1909 74817 1943 74851
rect 2053 74817 2087 74851
rect 2145 74817 2179 74851
rect 2329 74817 2363 74851
rect 3013 74817 3047 74851
rect 3433 74817 3467 74851
rect 1777 74681 1811 74715
rect 2881 74613 2915 74647
rect 2237 74341 2271 74375
rect 1409 74205 1443 74239
rect 2369 74205 2403 74239
rect 2513 74205 2547 74239
rect 2789 74205 2823 74239
rect 3985 74205 4019 74239
rect 10149 74205 10183 74239
rect 2605 74137 2639 74171
rect 1593 74069 1627 74103
rect 3801 74069 3835 74103
rect 9965 74069 9999 74103
rect 2513 73797 2547 73831
rect 2605 73797 2639 73831
rect 1409 73729 1443 73763
rect 2369 73729 2403 73763
rect 2789 73729 2823 73763
rect 1593 73593 1627 73627
rect 2237 73525 2271 73559
rect 2237 73253 2271 73287
rect 1409 73117 1443 73151
rect 2369 73117 2403 73151
rect 2789 73117 2823 73151
rect 10149 73117 10183 73151
rect 2513 73049 2547 73083
rect 2605 73049 2639 73083
rect 1593 72981 1627 73015
rect 9965 72981 9999 73015
rect 1409 72641 1443 72675
rect 2053 72641 2087 72675
rect 1593 72437 1627 72471
rect 2237 72437 2271 72471
rect 2237 72165 2271 72199
rect 1409 72029 1443 72063
rect 2369 72029 2403 72063
rect 2789 72029 2823 72063
rect 10149 72029 10183 72063
rect 2513 71961 2547 71995
rect 2605 71961 2639 71995
rect 1593 71893 1627 71927
rect 9965 71893 9999 71927
rect 2513 71621 2547 71655
rect 2605 71621 2639 71655
rect 1409 71553 1443 71587
rect 2369 71553 2403 71587
rect 2789 71553 2823 71587
rect 1593 71349 1627 71383
rect 2237 71349 2271 71383
rect 1961 71077 1995 71111
rect 1409 70941 1443 70975
rect 1829 70941 1863 70975
rect 2697 70941 2731 70975
rect 10149 70941 10183 70975
rect 1593 70873 1627 70907
rect 1685 70873 1719 70907
rect 2513 70805 2547 70839
rect 9965 70805 9999 70839
rect 2881 70533 2915 70567
rect 2697 70465 2731 70499
rect 2973 70465 3007 70499
rect 3070 70465 3104 70499
rect 1409 70397 1443 70431
rect 1685 70397 1719 70431
rect 3249 70329 3283 70363
rect 9965 70057 9999 70091
rect 1685 69921 1719 69955
rect 1409 69853 1443 69887
rect 2881 69853 2915 69887
rect 10149 69853 10183 69887
rect 2697 69717 2731 69751
rect 3157 69377 3191 69411
rect 4445 69377 4479 69411
rect 1409 69309 1443 69343
rect 1685 69309 1719 69343
rect 2881 69309 2915 69343
rect 4169 69309 4203 69343
rect 3893 68901 3927 68935
rect 1409 68765 1443 68799
rect 1685 68765 1719 68799
rect 4025 68765 4059 68799
rect 4445 68765 4479 68799
rect 10149 68765 10183 68799
rect 4169 68697 4203 68731
rect 4261 68697 4295 68731
rect 9965 68629 9999 68663
rect 4261 68357 4295 68391
rect 1680 68289 1714 68323
rect 1776 68289 1810 68323
rect 1869 68289 1903 68323
rect 2053 68289 2087 68323
rect 2605 68289 2639 68323
rect 2881 68289 2915 68323
rect 4117 68289 4151 68323
rect 4353 68289 4387 68323
rect 4537 68289 4571 68323
rect 1501 68085 1535 68119
rect 3985 68085 4019 68119
rect 9965 67881 9999 67915
rect 2881 67745 2915 67779
rect 3157 67745 3191 67779
rect 10149 67677 10183 67711
rect 1685 67609 1719 67643
rect 1869 67609 1903 67643
rect 1409 67201 1443 67235
rect 1685 67133 1719 67167
rect 1961 66521 1995 66555
rect 2697 66521 2731 66555
rect 1869 66453 1903 66487
rect 2605 66453 2639 66487
rect 9965 66249 9999 66283
rect 1961 66113 1995 66147
rect 2881 66113 2915 66147
rect 10149 66113 10183 66147
rect 1777 65977 1811 66011
rect 3065 65909 3099 65943
rect 2789 65501 2823 65535
rect 1777 65433 1811 65467
rect 1961 65433 1995 65467
rect 2605 65365 2639 65399
rect 1685 65025 1719 65059
rect 2789 65025 2823 65059
rect 10149 65025 10183 65059
rect 1501 64889 1535 64923
rect 2973 64821 3007 64855
rect 9965 64821 9999 64855
rect 2145 64549 2179 64583
rect 2324 64413 2358 64447
rect 2421 64413 2455 64447
rect 2697 64413 2731 64447
rect 3801 64413 3835 64447
rect 2513 64345 2547 64379
rect 3985 64277 4019 64311
rect 9965 64073 9999 64107
rect 2513 64005 2547 64039
rect 2605 64005 2639 64039
rect 1685 63937 1719 63971
rect 2369 63937 2403 63971
rect 2789 63937 2823 63971
rect 10149 63937 10183 63971
rect 1501 63733 1535 63767
rect 2237 63733 2271 63767
rect 2421 63393 2455 63427
rect 1685 63325 1719 63359
rect 3801 63325 3835 63359
rect 1501 63189 1535 63223
rect 2651 63189 2685 63223
rect 3985 63189 4019 63223
rect 9965 62985 9999 63019
rect 1961 62917 1995 62951
rect 2053 62917 2087 62951
rect 1864 62849 1898 62883
rect 2237 62849 2271 62883
rect 2973 62849 3007 62883
rect 10149 62849 10183 62883
rect 2697 62781 2731 62815
rect 1685 62645 1719 62679
rect 2237 62373 2271 62407
rect 1685 62237 1719 62271
rect 2369 62237 2403 62271
rect 2789 62237 2823 62271
rect 2513 62169 2547 62203
rect 2605 62169 2639 62203
rect 1501 62101 1535 62135
rect 2513 61829 2547 61863
rect 1685 61761 1719 61795
rect 2369 61761 2403 61795
rect 2605 61761 2639 61795
rect 2789 61761 2823 61795
rect 10149 61761 10183 61795
rect 9965 61625 9999 61659
rect 1501 61557 1535 61591
rect 2237 61557 2271 61591
rect 2237 61353 2271 61387
rect 1685 61149 1719 61183
rect 2421 61149 2455 61183
rect 1501 61013 1535 61047
rect 949 60809 983 60843
rect 9965 60809 9999 60843
rect 765 53533 799 53567
rect 857 52309 891 52343
rect 1685 60673 1719 60707
rect 10149 60673 10183 60707
rect 1501 60469 1535 60503
rect 1685 60061 1719 60095
rect 1501 59925 1535 59959
rect 1685 59585 1719 59619
rect 2421 59585 2455 59619
rect 10149 59585 10183 59619
rect 2237 59449 2271 59483
rect 1501 59381 1535 59415
rect 9965 59381 9999 59415
rect 1409 59109 1443 59143
rect 1593 58973 1627 59007
rect 1685 58973 1719 59007
rect 1961 58973 1995 59007
rect 2697 58973 2731 59007
rect 1777 58905 1811 58939
rect 2513 58837 2547 58871
rect 1685 58565 1719 58599
rect 1593 58497 1627 58531
rect 1777 58497 1811 58531
rect 1961 58497 1995 58531
rect 2697 58497 2731 58531
rect 10149 58497 10183 58531
rect 9965 58361 9999 58395
rect 1409 58293 1443 58327
rect 2513 58293 2547 58327
rect 1409 57885 1443 57919
rect 1685 57885 1719 57919
rect 1777 57885 1811 57919
rect 2421 57885 2455 57919
rect 2697 57885 2731 57919
rect 1593 57817 1627 57851
rect 1961 57749 1995 57783
rect 1593 57477 1627 57511
rect 1409 57409 1443 57443
rect 1685 57409 1719 57443
rect 1777 57409 1811 57443
rect 2697 57409 2731 57443
rect 3709 57409 3743 57443
rect 10149 57409 10183 57443
rect 2421 57341 2455 57375
rect 3893 57273 3927 57307
rect 1961 57205 1995 57239
rect 9965 57205 9999 57239
rect 1593 56797 1627 56831
rect 1961 56797 1995 56831
rect 2697 56797 2731 56831
rect 1685 56729 1719 56763
rect 1777 56729 1811 56763
rect 1409 56661 1443 56695
rect 2513 56661 2547 56695
rect 3065 56457 3099 56491
rect 9965 56457 9999 56491
rect 1685 56321 1719 56355
rect 2145 56321 2179 56355
rect 2973 56321 3007 56355
rect 10149 56321 10183 56355
rect 2329 56185 2363 56219
rect 1501 56117 1535 56151
rect 1685 55709 1719 55743
rect 1501 55573 1535 55607
rect 9965 55369 9999 55403
rect 1685 55233 1719 55267
rect 2421 55233 2455 55267
rect 10149 55233 10183 55267
rect 1501 55029 1535 55063
rect 2237 55029 2271 55063
rect 1685 54621 1719 54655
rect 1501 54485 1535 54519
rect 1685 54145 1719 54179
rect 2421 54145 2455 54179
rect 10149 54145 10183 54179
rect 2237 54009 2271 54043
rect 1501 53941 1535 53975
rect 9965 53941 9999 53975
rect 2881 53737 2915 53771
rect 1685 53533 1719 53567
rect 2145 53533 2179 53567
rect 2881 53533 2915 53567
rect 3065 53533 3099 53567
rect 1501 53397 1535 53431
rect 2329 53397 2363 53431
rect 3249 53193 3283 53227
rect 1593 53125 1627 53159
rect 1409 53057 1443 53091
rect 1685 53057 1719 53091
rect 1777 53057 1811 53091
rect 2697 53057 2731 53091
rect 3157 53057 3191 53091
rect 3341 53057 3375 53091
rect 10149 53057 10183 53091
rect 1961 52853 1995 52887
rect 2513 52853 2547 52887
rect 9965 52853 9999 52887
rect 3801 52649 3835 52683
rect 2789 52581 2823 52615
rect 1593 52445 1627 52479
rect 1777 52445 1811 52479
rect 1961 52445 1995 52479
rect 2605 52445 2639 52479
rect 3801 52445 3835 52479
rect 3985 52445 4019 52479
rect 1685 52377 1719 52411
rect 1409 52309 1443 52343
rect 949 52105 983 52139
rect 2513 51969 2547 52003
rect 10149 51969 10183 52003
rect 2237 51901 2271 51935
rect 2973 51901 3007 51935
rect 3249 51901 3283 51935
rect 857 51017 891 51051
rect 949 51765 983 51799
rect 9965 51765 9999 51799
rect 1409 51357 1443 51391
rect 1593 51357 1627 51391
rect 1777 51357 1811 51391
rect 2605 51357 2639 51391
rect 2973 51357 3007 51391
rect 3801 51357 3835 51391
rect 1685 51289 1719 51323
rect 2697 51289 2731 51323
rect 2789 51289 2823 51323
rect 1961 51221 1995 51255
rect 2421 51221 2455 51255
rect 3985 51221 4019 51255
rect 3433 51017 3467 51051
rect 9965 51017 9999 51051
rect 1961 50881 1995 50915
rect 3274 50881 3308 50915
rect 3985 50881 4019 50915
rect 4169 50881 4203 50915
rect 10149 50881 10183 50915
rect 765 49317 799 49351
rect 2237 50813 2271 50847
rect 213 46733 247 46767
rect 213 46053 247 46087
rect 3985 50677 4019 50711
rect 3801 50337 3835 50371
rect 4077 50337 4111 50371
rect 1593 50269 1627 50303
rect 1961 50269 1995 50303
rect 2697 50269 2731 50303
rect 1685 50201 1719 50235
rect 1777 50201 1811 50235
rect 1409 50133 1443 50167
rect 2513 50133 2547 50167
rect 1501 49929 1535 49963
rect 2973 49929 3007 49963
rect 9965 49929 9999 49963
rect 3617 49861 3651 49895
rect 1685 49793 1719 49827
rect 2421 49793 2455 49827
rect 2881 49793 2915 49827
rect 3065 49793 3099 49827
rect 3525 49793 3559 49827
rect 3709 49793 3743 49827
rect 10149 49793 10183 49827
rect 2237 49589 2271 49623
rect 2605 49385 2639 49419
rect 3065 49317 3099 49351
rect 3801 49249 3835 49283
rect 1685 49181 1719 49215
rect 2421 49181 2455 49215
rect 2605 49181 2639 49215
rect 3065 49181 3099 49215
rect 3249 49181 3283 49215
rect 4077 49181 4111 49215
rect 1501 49045 1535 49079
rect 1685 48705 1719 48739
rect 2421 48705 2455 48739
rect 10149 48705 10183 48739
rect 2237 48569 2271 48603
rect 1501 48501 1535 48535
rect 9965 48501 9999 48535
rect 10977 48501 11011 48535
rect 949 48297 983 48331
rect 2513 48229 2547 48263
rect 1685 48093 1719 48127
rect 2513 48093 2547 48127
rect 2697 48093 2731 48127
rect 1501 47957 1535 47991
rect 2973 47685 3007 47719
rect 1685 47617 1719 47651
rect 2421 47617 2455 47651
rect 2881 47617 2915 47651
rect 3065 47617 3099 47651
rect 10149 47617 10183 47651
rect 1501 47413 1535 47447
rect 2237 47413 2271 47447
rect 9965 47413 9999 47447
rect 2513 47209 2547 47243
rect 3801 47209 3835 47243
rect 1685 47005 1719 47039
rect 2513 47005 2547 47039
rect 2697 47005 2731 47039
rect 3801 47005 3835 47039
rect 3985 47005 4019 47039
rect 1501 46869 1535 46903
rect 3709 46665 3743 46699
rect 1685 46529 1719 46563
rect 2421 46529 2455 46563
rect 2881 46529 2915 46563
rect 3617 46529 3651 46563
rect 3801 46529 3835 46563
rect 10149 46529 10183 46563
rect 3065 46393 3099 46427
rect 1501 46325 1535 46359
rect 2237 46325 2271 46359
rect 9965 46325 9999 46359
rect 2421 45985 2455 46019
rect 1685 45917 1719 45951
rect 2697 45917 2731 45951
rect 1501 45781 1535 45815
rect 2697 45441 2731 45475
rect 10149 45441 10183 45475
rect 2421 45373 2455 45407
rect 9965 45237 9999 45271
rect 1593 44829 1627 44863
rect 1961 44829 1995 44863
rect 2697 44829 2731 44863
rect 949 44761 983 44795
rect 1685 44761 1719 44795
rect 1777 44761 1811 44795
rect 1409 44693 1443 44727
rect 2513 44693 2547 44727
rect 11069 47413 11103 47447
rect 11069 44761 11103 44795
rect 10977 44489 11011 44523
rect 1685 44421 1719 44455
rect 2697 44421 2731 44455
rect 2789 44421 2823 44455
rect 1593 44353 1627 44387
rect 1777 44353 1811 44387
rect 1961 44353 1995 44387
rect 2605 44353 2639 44387
rect 2973 44353 3007 44387
rect 10149 44353 10183 44387
rect 1409 44149 1443 44183
rect 2421 44149 2455 44183
rect 9965 44149 9999 44183
rect 1593 43741 1627 43775
rect 1685 43741 1719 43775
rect 1961 43741 1995 43775
rect 2421 43741 2455 43775
rect 3801 43741 3835 43775
rect 1777 43673 1811 43707
rect 1409 43605 1443 43639
rect 2605 43605 2639 43639
rect 3985 43605 4019 43639
rect 1777 43333 1811 43367
rect 1593 43265 1627 43299
rect 1685 43265 1719 43299
rect 1961 43265 1995 43299
rect 2697 43265 2731 43299
rect 9873 43265 9907 43299
rect 857 42245 891 42279
rect 949 43061 983 43095
rect 1409 43061 1443 43095
rect 2513 43061 2547 43095
rect 10057 43061 10091 43095
rect 857 42109 891 42143
rect 4721 42857 4755 42891
rect 1685 42653 1719 42687
rect 2421 42653 2455 42687
rect 4537 42653 4571 42687
rect 4721 42653 4755 42687
rect 1501 42517 1535 42551
rect 2237 42517 2271 42551
rect 1685 42177 1719 42211
rect 4537 42177 4571 42211
rect 4721 42177 4755 42211
rect 9873 42177 9907 42211
rect 4629 42109 4663 42143
rect 1501 41973 1535 42007
rect 10057 41973 10091 42007
rect 1685 41565 1719 41599
rect 1501 41429 1535 41463
rect 1685 41089 1719 41123
rect 4537 41089 4571 41123
rect 4721 41089 4755 41123
rect 9873 41089 9907 41123
rect 1501 40885 1535 40919
rect 4721 40885 4755 40919
rect 10057 40885 10091 40919
rect 1685 40477 1719 40511
rect 1501 40341 1535 40375
rect 2605 40137 2639 40171
rect 1685 40001 1719 40035
rect 2513 40001 2547 40035
rect 2697 40001 2731 40035
rect 1501 39797 1535 39831
rect 2421 39525 2455 39559
rect 1685 39389 1719 39423
rect 2513 39389 2547 39423
rect 2697 39389 2731 39423
rect 9873 39389 9907 39423
rect 1501 39253 1535 39287
rect 10057 39253 10091 39287
rect 2329 38981 2363 39015
rect 1685 38913 1719 38947
rect 2513 38913 2547 38947
rect 2605 38913 2639 38947
rect 4261 38913 4295 38947
rect 4445 38913 4479 38947
rect 1501 38777 1535 38811
rect 4445 38709 4479 38743
rect 2421 38437 2455 38471
rect 1685 38301 1719 38335
rect 2513 38301 2547 38335
rect 2605 38301 2639 38335
rect 4261 38301 4295 38335
rect 4445 38301 4479 38335
rect 9873 38301 9907 38335
rect 1501 38165 1535 38199
rect 4353 38165 4387 38199
rect 10057 38165 10091 38199
rect 1501 37961 1535 37995
rect 2513 37961 2547 37995
rect 1685 37825 1719 37859
rect 2237 37825 2271 37859
rect 2513 37825 2547 37859
rect 3065 37825 3099 37859
rect 4169 37825 4203 37859
rect 4353 37825 4387 37859
rect 3249 37621 3283 37655
rect 4353 37621 4387 37655
rect 1409 37213 1443 37247
rect 2145 37213 2179 37247
rect 2973 37213 3007 37247
rect 3065 37213 3099 37247
rect 9873 37213 9907 37247
rect 1593 37077 1627 37111
rect 2329 37077 2363 37111
rect 10057 37077 10091 37111
rect 2237 36873 2271 36907
rect 2881 36873 2915 36907
rect 949 36805 983 36839
rect 1685 36737 1719 36771
rect 2329 36737 2363 36771
rect 2789 36737 2823 36771
rect 4169 36737 4203 36771
rect 4353 36737 4387 36771
rect 1501 36533 1535 36567
rect 4353 36533 4387 36567
rect 2237 36329 2271 36363
rect 1409 36125 1443 36159
rect 2329 36125 2363 36159
rect 4169 36125 4203 36159
rect 4353 36125 4387 36159
rect 9873 36125 9907 36159
rect 857 36057 891 36091
rect 1593 35989 1627 36023
rect 4261 35989 4295 36023
rect 10057 35989 10091 36023
rect 2973 35785 3007 35819
rect 1685 35649 1719 35683
rect 2145 35649 2179 35683
rect 3157 35649 3191 35683
rect 2329 35513 2363 35547
rect 1501 35445 1535 35479
rect 4537 35105 4571 35139
rect 1409 35037 1443 35071
rect 4261 35037 4295 35071
rect 9873 35037 9907 35071
rect 1593 34901 1627 34935
rect 10057 34901 10091 34935
rect 2329 34697 2363 34731
rect 3249 34629 3283 34663
rect 1409 34561 1443 34595
rect 2513 34561 2547 34595
rect 3065 34561 3099 34595
rect 1593 34357 1627 34391
rect 3065 34153 3099 34187
rect 1409 33949 1443 33983
rect 2329 33949 2363 33983
rect 2513 33949 2547 33983
rect 3249 33949 3283 33983
rect 9873 33949 9907 33983
rect 1593 33813 1627 33847
rect 2513 33813 2547 33847
rect 10057 33813 10091 33847
rect 2513 33609 2547 33643
rect 3157 33609 3191 33643
rect 1777 33473 1811 33507
rect 2329 33473 2363 33507
rect 2513 33473 2547 33507
rect 3157 33473 3191 33507
rect 3433 33473 3467 33507
rect 4353 33473 4387 33507
rect 4537 33473 4571 33507
rect 1777 33269 1811 33303
rect 4537 33269 4571 33303
rect 3065 33065 3099 33099
rect 1593 32997 1627 33031
rect 2329 32997 2363 33031
rect 1409 32861 1443 32895
rect 2421 32861 2455 32895
rect 2605 32861 2639 32895
rect 3249 32861 3283 32895
rect 4353 32861 4387 32895
rect 4537 32861 4571 32895
rect 9873 32861 9907 32895
rect 4445 32725 4479 32759
rect 10057 32725 10091 32759
rect 1593 32521 1627 32555
rect 2237 32453 2271 32487
rect 3157 32453 3191 32487
rect 1409 32385 1443 32419
rect 2421 32385 2455 32419
rect 2513 32385 2547 32419
rect 4629 32385 4663 32419
rect 3341 32317 3375 32351
rect 4353 32317 4387 32351
rect 1961 31977 1995 32011
rect 2513 31977 2547 32011
rect 4537 31841 4571 31875
rect 2053 31773 2087 31807
rect 2697 31773 2731 31807
rect 4445 31773 4479 31807
rect 4629 31773 4663 31807
rect 9873 31773 9907 31807
rect 10057 31637 10091 31671
rect 2421 31433 2455 31467
rect 1777 31365 1811 31399
rect 1869 31297 1903 31331
rect 2329 31297 2363 31331
rect 4445 31297 4479 31331
rect 4629 31297 4663 31331
rect 4629 31093 4663 31127
rect 1777 30889 1811 30923
rect 2329 30889 2363 30923
rect 3801 30889 3835 30923
rect 2973 30821 3007 30855
rect 1869 30685 1903 30719
rect 2513 30685 2547 30719
rect 3157 30685 3191 30719
rect 3985 30685 4019 30719
rect 4445 30685 4479 30719
rect 4629 30685 4663 30719
rect 9873 30685 9907 30719
rect 4537 30549 4571 30583
rect 10057 30549 10091 30583
rect 2513 30345 2547 30379
rect 1869 30209 1903 30243
rect 2329 30209 2363 30243
rect 1777 30141 1811 30175
rect 2421 29801 2455 29835
rect 3065 29801 3099 29835
rect 1869 29665 1903 29699
rect 1961 29597 1995 29631
rect 2605 29597 2639 29631
rect 3249 29597 3283 29631
rect 9873 29597 9907 29631
rect 10057 29461 10091 29495
rect 2145 29257 2179 29291
rect 2697 29257 2731 29291
rect 3341 29257 3375 29291
rect 1961 29121 1995 29155
rect 2145 29121 2179 29155
rect 2881 29121 2915 29155
rect 3525 29121 3559 29155
rect 2789 28645 2823 28679
rect 1869 28577 1903 28611
rect 2053 28509 2087 28543
rect 2145 28509 2179 28543
rect 2881 28509 2915 28543
rect 3065 28509 3099 28543
rect 3801 28509 3835 28543
rect 3985 28509 4019 28543
rect 9873 28509 9907 28543
rect 3893 28373 3927 28407
rect 10057 28373 10091 28407
rect 2973 28169 3007 28203
rect 2237 28101 2271 28135
rect 1869 28033 1903 28067
rect 2145 28033 2179 28067
rect 2881 28033 2915 28067
rect 3065 28033 3099 28067
rect 3985 28033 4019 28067
rect 4261 27965 4295 27999
rect 2881 27625 2915 27659
rect 1501 27557 1535 27591
rect 2053 27557 2087 27591
rect 1593 27421 1627 27455
rect 2237 27421 2271 27455
rect 2973 27421 3007 27455
rect 3801 27421 3835 27455
rect 3985 27421 4019 27455
rect 9873 27421 9907 27455
rect 3893 27285 3927 27319
rect 10057 27285 10091 27319
rect 2697 27081 2731 27115
rect 2145 27013 2179 27047
rect 1593 26945 1627 26979
rect 2053 26945 2087 26979
rect 2881 26945 2915 26979
rect 3617 26945 3651 26979
rect 3801 26945 3835 26979
rect 1501 26877 1535 26911
rect 3801 26741 3835 26775
rect 2237 26537 2271 26571
rect 3985 26537 4019 26571
rect 1501 26469 1535 26503
rect 4629 26469 4663 26503
rect 2881 26401 2915 26435
rect 1593 26333 1627 26367
rect 2053 26333 2087 26367
rect 3801 26333 3835 26367
rect 3985 26333 4019 26367
rect 4445 26333 4479 26367
rect 4629 26333 4663 26367
rect 9873 26333 9907 26367
rect 3157 26265 3191 26299
rect 10057 26197 10091 26231
rect 1501 25993 1535 26027
rect 2053 25993 2087 26027
rect 1593 25857 1627 25891
rect 2237 25857 2271 25891
rect 2053 25449 2087 25483
rect 2697 25381 2731 25415
rect 1409 25245 1443 25279
rect 2237 25245 2271 25279
rect 2881 25245 2915 25279
rect 9873 25245 9907 25279
rect 1593 25109 1627 25143
rect 10057 25109 10091 25143
rect 1409 24769 1443 24803
rect 3249 24769 3283 24803
rect 3341 24769 3375 24803
rect 4077 24769 4111 24803
rect 1593 24565 1627 24599
rect 4353 24565 4387 24599
rect 2697 24293 2731 24327
rect 4445 24293 4479 24327
rect 1593 24157 1627 24191
rect 2053 24157 2087 24191
rect 2881 24157 2915 24191
rect 4261 24157 4295 24191
rect 9873 24157 9907 24191
rect 1501 24021 1535 24055
rect 2145 24021 2179 24055
rect 10057 24021 10091 24055
rect 3065 23817 3099 23851
rect 2053 23681 2087 23715
rect 2237 23681 2271 23715
rect 2973 23681 3007 23715
rect 3157 23681 3191 23715
rect 3801 23681 3835 23715
rect 2237 23545 2271 23579
rect 3617 23477 3651 23511
rect 3065 23273 3099 23307
rect 2053 23137 2087 23171
rect 1409 23069 1443 23103
rect 2237 23069 2271 23103
rect 2421 23069 2455 23103
rect 4077 23069 4111 23103
rect 4261 23069 4295 23103
rect 4721 23069 4755 23103
rect 4905 23069 4939 23103
rect 9873 23069 9907 23103
rect 1501 23001 1535 23035
rect 2973 23001 3007 23035
rect 4169 22933 4203 22967
rect 4813 22933 4847 22967
rect 10057 22933 10091 22967
rect 2145 22729 2179 22763
rect 3157 22729 3191 22763
rect 1409 22593 1443 22627
rect 2053 22593 2087 22627
rect 2329 22593 2363 22627
rect 2973 22593 3007 22627
rect 3249 22593 3283 22627
rect 4537 22593 4571 22627
rect 1501 22525 1535 22559
rect 4261 22525 4295 22559
rect 2881 22185 2915 22219
rect 1593 21981 1627 22015
rect 2053 21981 2087 22015
rect 2973 21981 3007 22015
rect 4077 21981 4111 22015
rect 4261 21981 4295 22015
rect 9873 21981 9907 22015
rect 1501 21845 1535 21879
rect 2237 21845 2271 21879
rect 4169 21845 4203 21879
rect 10057 21845 10091 21879
rect 1593 21641 1627 21675
rect 1409 21505 1443 21539
rect 2237 21505 2271 21539
rect 2881 21505 2915 21539
rect 3341 21505 3375 21539
rect 4077 21505 4111 21539
rect 4261 21505 4295 21539
rect 4721 21505 4755 21539
rect 4905 21505 4939 21539
rect 4261 21369 4295 21403
rect 10977 21369 11011 21403
rect 2053 21301 2087 21335
rect 2697 21301 2731 21335
rect 3525 21301 3559 21335
rect 4905 21301 4939 21335
rect 4445 20961 4479 20995
rect 1409 20893 1443 20927
rect 2237 20893 2271 20927
rect 3065 20893 3099 20927
rect 4721 20893 4755 20927
rect 9873 20893 9907 20927
rect 1593 20757 1627 20791
rect 2053 20757 2087 20791
rect 2881 20757 2915 20791
rect 10057 20757 10091 20791
rect 2145 20485 2179 20519
rect 1409 20417 1443 20451
rect 2237 20417 2271 20451
rect 2697 20417 2731 20451
rect 3525 20417 3559 20451
rect 2789 20281 2823 20315
rect 1593 20213 1627 20247
rect 3341 20213 3375 20247
rect 2421 19941 2455 19975
rect 1869 19805 1903 19839
rect 2513 19805 2547 19839
rect 2697 19805 2731 19839
rect 3801 19805 3835 19839
rect 9873 19805 9907 19839
rect 1777 19737 1811 19771
rect 3893 19669 3927 19703
rect 10057 19669 10091 19703
rect 1777 19465 1811 19499
rect 2973 19465 3007 19499
rect 3801 19465 3835 19499
rect 1685 19329 1719 19363
rect 1869 19329 1903 19363
rect 2513 19329 2547 19363
rect 3065 19329 3099 19363
rect 3617 19329 3651 19363
rect 3893 19329 3927 19363
rect 1777 18921 1811 18955
rect 1869 18717 1903 18751
rect 2513 18717 2547 18751
rect 3065 18717 3099 18751
rect 3985 18717 4019 18751
rect 9873 18717 9907 18751
rect 10977 18717 11011 18751
rect 2973 18581 3007 18615
rect 3801 18581 3835 18615
rect 10057 18581 10091 18615
rect 2145 18377 2179 18411
rect 1409 18241 1443 18275
rect 2053 18241 2087 18275
rect 2881 18241 2915 18275
rect 3525 18241 3559 18275
rect 4353 18241 4387 18275
rect 4537 18241 4571 18275
rect 4997 18241 5031 18275
rect 5181 18241 5215 18275
rect 2789 18105 2823 18139
rect 4537 18105 4571 18139
rect 1593 18037 1627 18071
rect 3341 18037 3375 18071
rect 5181 18037 5215 18071
rect 2145 17833 2179 17867
rect 1409 17629 1443 17663
rect 2053 17629 2087 17663
rect 2881 17629 2915 17663
rect 4353 17629 4387 17663
rect 4537 17629 4571 17663
rect 4997 17629 5031 17663
rect 5181 17629 5215 17663
rect 9873 17629 9907 17663
rect 10977 17561 11011 17595
rect 1593 17493 1627 17527
rect 2697 17493 2731 17527
rect 4445 17493 4479 17527
rect 5089 17493 5123 17527
rect 10057 17493 10091 17527
rect 2145 17289 2179 17323
rect 1409 17153 1443 17187
rect 2237 17153 2271 17187
rect 4353 17153 4387 17187
rect 4537 17153 4571 17187
rect 1593 16949 1627 16983
rect 4537 16949 4571 16983
rect 1961 16745 1995 16779
rect 1501 16609 1535 16643
rect 1593 16541 1627 16575
rect 1961 16541 1995 16575
rect 9873 16541 9907 16575
rect 2145 16405 2179 16439
rect 10057 16405 10091 16439
rect 1409 16065 1443 16099
rect 2237 16065 2271 16099
rect 1593 15929 1627 15963
rect 2053 15861 2087 15895
rect 1409 15453 1443 15487
rect 2237 15453 2271 15487
rect 9873 15453 9907 15487
rect 1593 15317 1627 15351
rect 2053 15317 2087 15351
rect 10057 15317 10091 15351
rect 1593 15045 1627 15079
rect 1409 14977 1443 15011
rect 1777 14773 1811 14807
rect 1869 14569 1903 14603
rect 1409 14501 1443 14535
rect 1777 14433 1811 14467
rect 1593 14365 1627 14399
rect 1869 14365 1903 14399
rect 2329 14365 2363 14399
rect 9873 14365 9907 14399
rect 10977 14365 11011 14399
rect 11069 17289 11103 17323
rect 2513 14229 2547 14263
rect 10057 14229 10091 14263
rect 1593 14025 1627 14059
rect 2053 14025 2087 14059
rect 1409 13889 1443 13923
rect 2237 13889 2271 13923
rect 1409 13277 1443 13311
rect 1593 13141 1627 13175
rect 1409 12801 1443 12835
rect 2237 12801 2271 12835
rect 9873 12801 9907 12835
rect 11069 12801 11103 12835
rect 10057 12665 10091 12699
rect 1593 12597 1627 12631
rect 2053 12597 2087 12631
rect 1593 12189 1627 12223
rect 2237 12189 2271 12223
rect 1409 12121 1443 12155
rect 1777 12053 1811 12087
rect 2329 12053 2363 12087
rect 1869 11849 1903 11883
rect 2697 11781 2731 11815
rect 1409 11713 1443 11747
rect 1685 11713 1719 11747
rect 2329 11713 2363 11747
rect 3985 11713 4019 11747
rect 4169 11713 4203 11747
rect 9873 11713 9907 11747
rect 1593 11645 1627 11679
rect 2421 11645 2455 11679
rect 2697 11577 2731 11611
rect 4169 11577 4203 11611
rect 10057 11577 10091 11611
rect 1685 11509 1719 11543
rect 2513 11509 2547 11543
rect 2697 11169 2731 11203
rect 1409 11101 1443 11135
rect 2145 11101 2179 11135
rect 2237 11101 2271 11135
rect 2421 11101 2455 11135
rect 3985 11101 4019 11135
rect 4169 11101 4203 11135
rect 4077 11033 4111 11067
rect 1593 10965 1627 10999
rect 2697 10761 2731 10795
rect 2053 10625 2087 10659
rect 2237 10625 2271 10659
rect 2513 10625 2547 10659
rect 4353 10625 4387 10659
rect 9873 10625 9907 10659
rect 4629 10557 4663 10591
rect 10057 10489 10091 10523
rect 1593 10217 1627 10251
rect 1961 10217 1995 10251
rect 1685 10081 1719 10115
rect 1409 10013 1443 10047
rect 3985 10013 4019 10047
rect 4169 10013 4203 10047
rect 4077 9877 4111 9911
rect 3985 9537 4019 9571
rect 4169 9537 4203 9571
rect 4813 9537 4847 9571
rect 9873 9537 9907 9571
rect 5089 9469 5123 9503
rect 10057 9401 10091 9435
rect 4169 9333 4203 9367
rect 9873 8449 9907 8483
rect 10057 8313 10091 8347
rect 3893 7837 3927 7871
rect 4077 7837 4111 7871
rect 3985 7701 4019 7735
rect 9873 7361 9907 7395
rect 10057 7225 10091 7259
rect 4629 6749 4663 6783
rect 4813 6749 4847 6783
rect 4721 6613 4755 6647
rect 2881 6409 2915 6443
rect 2237 6341 2271 6375
rect 2145 6273 2179 6307
rect 2789 6273 2823 6307
rect 4629 6273 4663 6307
rect 4813 6273 4847 6307
rect 9873 6273 9907 6307
rect 4813 6069 4847 6103
rect 10057 6069 10091 6103
rect 2237 5865 2271 5899
rect 3985 5865 4019 5899
rect 11069 5865 11103 5899
rect 1593 5797 1627 5831
rect 2881 5797 2915 5831
rect 3617 5797 3651 5831
rect 1409 5661 1443 5695
rect 2145 5661 2179 5695
rect 2789 5661 2823 5695
rect 3801 5661 3835 5695
rect 4629 5661 4663 5695
rect 4813 5661 4847 5695
rect 5261 5661 5295 5695
rect 5457 5661 5491 5695
rect 4721 5593 4755 5627
rect 10977 5593 11011 5627
rect 3617 5525 3651 5559
rect 5365 5525 5399 5559
rect 2237 5321 2271 5355
rect 2881 5321 2915 5355
rect 2145 5185 2179 5219
rect 2789 5185 2823 5219
rect 4629 5185 4663 5219
rect 4813 5185 4847 5219
rect 9873 5185 9907 5219
rect 4813 4981 4847 5015
rect 10057 4981 10091 5015
rect 1593 4777 1627 4811
rect 1409 4573 1443 4607
rect 1409 4097 1443 4131
rect 9873 4097 9907 4131
rect 1593 3961 1627 3995
rect 10057 3893 10091 3927
rect 1593 3689 1627 3723
rect 1409 3485 1443 3519
rect 9873 3485 9907 3519
rect 10057 3349 10091 3383
rect 1593 3145 1627 3179
rect 1409 3009 1443 3043
rect 9873 3009 9907 3043
rect 10977 3009 11011 3043
rect 10057 2805 10091 2839
rect 10977 2805 11011 2839
rect 1593 2601 1627 2635
rect 2237 2601 2271 2635
rect 2881 2601 2915 2635
rect 1409 2397 1443 2431
rect 2053 2397 2087 2431
rect 2697 2397 2731 2431
rect 9873 2397 9907 2431
rect 10057 2261 10091 2295
rect 11069 2397 11103 2431
rect 10977 629 11011 663
<< metal1 >>
rect 10962 78248 10968 78260
rect 10923 78220 10968 78248
rect 10962 78208 10968 78220
rect 11020 78208 11026 78260
rect 1104 77818 10856 77840
rect 1104 77766 2582 77818
rect 2634 77766 2646 77818
rect 2698 77766 2710 77818
rect 2762 77766 2774 77818
rect 2826 77766 2838 77818
rect 2890 77766 5845 77818
rect 5897 77766 5909 77818
rect 5961 77766 5973 77818
rect 6025 77766 6037 77818
rect 6089 77766 6101 77818
rect 6153 77766 9109 77818
rect 9161 77766 9173 77818
rect 9225 77766 9237 77818
rect 9289 77766 9301 77818
rect 9353 77766 9365 77818
rect 9417 77766 10856 77818
rect 1104 77744 10856 77766
rect 1397 77503 1455 77509
rect 1397 77469 1409 77503
rect 1443 77500 1455 77503
rect 1486 77500 1492 77512
rect 1443 77472 1492 77500
rect 1443 77469 1455 77472
rect 1397 77463 1455 77469
rect 1486 77460 1492 77472
rect 1544 77460 1550 77512
rect 2038 77500 2044 77512
rect 1999 77472 2044 77500
rect 2038 77460 2044 77472
rect 2096 77460 2102 77512
rect 2866 77500 2872 77512
rect 2827 77472 2872 77500
rect 2866 77460 2872 77472
rect 2924 77460 2930 77512
rect 3970 77500 3976 77512
rect 3931 77472 3976 77500
rect 3970 77460 3976 77472
rect 4028 77460 4034 77512
rect 9490 77500 9496 77512
rect 9451 77472 9496 77500
rect 9490 77460 9496 77472
rect 9548 77460 9554 77512
rect 10134 77500 10140 77512
rect 10095 77472 10140 77500
rect 10134 77460 10140 77472
rect 10192 77460 10198 77512
rect 1578 77364 1584 77376
rect 1539 77336 1584 77364
rect 1578 77324 1584 77336
rect 1636 77324 1642 77376
rect 2130 77324 2136 77376
rect 2188 77364 2194 77376
rect 2225 77367 2283 77373
rect 2225 77364 2237 77367
rect 2188 77336 2237 77364
rect 2188 77324 2194 77336
rect 2225 77333 2237 77336
rect 2271 77333 2283 77367
rect 2225 77327 2283 77333
rect 2406 77324 2412 77376
rect 2464 77364 2470 77376
rect 2685 77367 2743 77373
rect 2685 77364 2697 77367
rect 2464 77336 2697 77364
rect 2464 77324 2470 77336
rect 2685 77333 2697 77336
rect 2731 77333 2743 77367
rect 2685 77327 2743 77333
rect 2866 77324 2872 77376
rect 2924 77364 2930 77376
rect 3789 77367 3847 77373
rect 3789 77364 3801 77367
rect 2924 77336 3801 77364
rect 2924 77324 2930 77336
rect 3789 77333 3801 77336
rect 3835 77333 3847 77367
rect 3789 77327 3847 77333
rect 5534 77324 5540 77376
rect 5592 77364 5598 77376
rect 9309 77367 9367 77373
rect 9309 77364 9321 77367
rect 5592 77336 9321 77364
rect 5592 77324 5598 77336
rect 9309 77333 9321 77336
rect 9355 77333 9367 77367
rect 9309 77327 9367 77333
rect 9674 77324 9680 77376
rect 9732 77364 9738 77376
rect 9953 77367 10011 77373
rect 9953 77364 9965 77367
rect 9732 77336 9965 77364
rect 9732 77324 9738 77336
rect 9953 77333 9965 77336
rect 9999 77333 10011 77367
rect 9953 77327 10011 77333
rect 1104 77274 10856 77296
rect 1104 77222 4213 77274
rect 4265 77222 4277 77274
rect 4329 77222 4341 77274
rect 4393 77222 4405 77274
rect 4457 77222 4469 77274
rect 4521 77222 7477 77274
rect 7529 77222 7541 77274
rect 7593 77222 7605 77274
rect 7657 77222 7669 77274
rect 7721 77222 7733 77274
rect 7785 77222 10856 77274
rect 1104 77200 10856 77222
rect 1394 77024 1400 77036
rect 1355 76996 1400 77024
rect 1394 76984 1400 76996
rect 1452 76984 1458 77036
rect 2038 77024 2044 77036
rect 1999 76996 2044 77024
rect 2038 76984 2044 76996
rect 2096 76984 2102 77036
rect 2869 77027 2927 77033
rect 2869 76993 2881 77027
rect 2915 77024 2927 77027
rect 2958 77024 2964 77036
rect 2915 76996 2964 77024
rect 2915 76993 2927 76996
rect 2869 76987 2927 76993
rect 2958 76984 2964 76996
rect 3016 76984 3022 77036
rect 10137 77027 10195 77033
rect 10137 76993 10149 77027
rect 10183 77024 10195 77027
rect 10965 77027 11023 77033
rect 10965 77024 10977 77027
rect 10183 76996 10977 77024
rect 10183 76993 10195 76996
rect 10137 76987 10195 76993
rect 10965 76993 10977 76996
rect 11011 76993 11023 77027
rect 10965 76987 11023 76993
rect 1581 76823 1639 76829
rect 1581 76789 1593 76823
rect 1627 76820 1639 76823
rect 1670 76820 1676 76832
rect 1627 76792 1676 76820
rect 1627 76789 1639 76792
rect 1581 76783 1639 76789
rect 1670 76780 1676 76792
rect 1728 76780 1734 76832
rect 2225 76823 2283 76829
rect 2225 76789 2237 76823
rect 2271 76820 2283 76823
rect 2314 76820 2320 76832
rect 2271 76792 2320 76820
rect 2271 76789 2283 76792
rect 2225 76783 2283 76789
rect 2314 76780 2320 76792
rect 2372 76780 2378 76832
rect 2498 76780 2504 76832
rect 2556 76820 2562 76832
rect 2685 76823 2743 76829
rect 2685 76820 2697 76823
rect 2556 76792 2697 76820
rect 2556 76780 2562 76792
rect 2685 76789 2697 76792
rect 2731 76789 2743 76823
rect 9950 76820 9956 76832
rect 9911 76792 9956 76820
rect 2685 76783 2743 76789
rect 9950 76780 9956 76792
rect 10008 76780 10014 76832
rect 1104 76730 10856 76752
rect 1104 76678 2582 76730
rect 2634 76678 2646 76730
rect 2698 76678 2710 76730
rect 2762 76678 2774 76730
rect 2826 76678 2838 76730
rect 2890 76678 5845 76730
rect 5897 76678 5909 76730
rect 5961 76678 5973 76730
rect 6025 76678 6037 76730
rect 6089 76678 6101 76730
rect 6153 76678 9109 76730
rect 9161 76678 9173 76730
rect 9225 76678 9237 76730
rect 9289 76678 9301 76730
rect 9353 76678 9365 76730
rect 9417 76678 10856 76730
rect 1104 76656 10856 76678
rect 3050 76480 3056 76492
rect 2240 76452 3056 76480
rect 1302 76372 1308 76424
rect 1360 76412 1366 76424
rect 2240 76421 2268 76452
rect 3050 76440 3056 76452
rect 3108 76440 3114 76492
rect 1397 76415 1455 76421
rect 1397 76412 1409 76415
rect 1360 76384 1409 76412
rect 1360 76372 1366 76384
rect 1397 76381 1409 76384
rect 1443 76381 1455 76415
rect 1397 76375 1455 76381
rect 2225 76415 2283 76421
rect 2225 76381 2237 76415
rect 2271 76381 2283 76415
rect 2225 76375 2283 76381
rect 2685 76415 2743 76421
rect 2685 76381 2697 76415
rect 2731 76412 2743 76415
rect 3142 76412 3148 76424
rect 2731 76384 3148 76412
rect 2731 76381 2743 76384
rect 2685 76375 2743 76381
rect 3142 76372 3148 76384
rect 3200 76372 3206 76424
rect 10134 76412 10140 76424
rect 10095 76384 10140 76412
rect 10134 76372 10140 76384
rect 10192 76372 10198 76424
rect 3510 76344 3516 76356
rect 1596 76316 3516 76344
rect 1596 76285 1624 76316
rect 3510 76304 3516 76316
rect 3568 76304 3574 76356
rect 1581 76279 1639 76285
rect 1581 76245 1593 76279
rect 1627 76245 1639 76279
rect 2038 76276 2044 76288
rect 1999 76248 2044 76276
rect 1581 76239 1639 76245
rect 2038 76236 2044 76248
rect 2096 76236 2102 76288
rect 2869 76279 2927 76285
rect 2869 76245 2881 76279
rect 2915 76276 2927 76279
rect 3142 76276 3148 76288
rect 2915 76248 3148 76276
rect 2915 76245 2927 76248
rect 2869 76239 2927 76245
rect 3142 76236 3148 76248
rect 3200 76236 3206 76288
rect 9766 76236 9772 76288
rect 9824 76276 9830 76288
rect 9953 76279 10011 76285
rect 9953 76276 9965 76279
rect 9824 76248 9965 76276
rect 9824 76236 9830 76248
rect 9953 76245 9965 76248
rect 9999 76245 10011 76279
rect 9953 76239 10011 76245
rect 1104 76186 10856 76208
rect 1104 76134 4213 76186
rect 4265 76134 4277 76186
rect 4329 76134 4341 76186
rect 4393 76134 4405 76186
rect 4457 76134 4469 76186
rect 4521 76134 7477 76186
rect 7529 76134 7541 76186
rect 7593 76134 7605 76186
rect 7657 76134 7669 76186
rect 7721 76134 7733 76186
rect 7785 76134 10856 76186
rect 1104 76112 10856 76134
rect 1581 76075 1639 76081
rect 1581 76041 1593 76075
rect 1627 76072 1639 76075
rect 1854 76072 1860 76084
rect 1627 76044 1860 76072
rect 1627 76041 1639 76044
rect 1581 76035 1639 76041
rect 1854 76032 1860 76044
rect 1912 76032 1918 76084
rect 1946 76032 1952 76084
rect 2004 76072 2010 76084
rect 2041 76075 2099 76081
rect 2041 76072 2053 76075
rect 2004 76044 2053 76072
rect 2004 76032 2010 76044
rect 2041 76041 2053 76044
rect 2087 76041 2099 76075
rect 2041 76035 2099 76041
rect 1394 75936 1400 75948
rect 1355 75908 1400 75936
rect 1394 75896 1400 75908
rect 1452 75896 1458 75948
rect 1486 75896 1492 75948
rect 1544 75936 1550 75948
rect 1670 75936 1676 75948
rect 1544 75908 1676 75936
rect 1544 75896 1550 75908
rect 1670 75896 1676 75908
rect 1728 75896 1734 75948
rect 2222 75936 2228 75948
rect 2183 75908 2228 75936
rect 2222 75896 2228 75908
rect 2280 75896 2286 75948
rect 1104 75642 10856 75664
rect 1104 75590 2582 75642
rect 2634 75590 2646 75642
rect 2698 75590 2710 75642
rect 2762 75590 2774 75642
rect 2826 75590 2838 75642
rect 2890 75590 5845 75642
rect 5897 75590 5909 75642
rect 5961 75590 5973 75642
rect 6025 75590 6037 75642
rect 6089 75590 6101 75642
rect 6153 75590 9109 75642
rect 9161 75590 9173 75642
rect 9225 75590 9237 75642
rect 9289 75590 9301 75642
rect 9353 75590 9365 75642
rect 9417 75590 10856 75642
rect 1104 75568 10856 75590
rect 1118 75420 1124 75472
rect 1176 75460 1182 75472
rect 1765 75463 1823 75469
rect 1765 75460 1777 75463
rect 1176 75432 1777 75460
rect 1176 75420 1182 75432
rect 1765 75429 1777 75432
rect 1811 75429 1823 75463
rect 1765 75423 1823 75429
rect 1944 75327 2002 75333
rect 1944 75293 1956 75327
rect 1990 75293 2002 75327
rect 1944 75287 2002 75293
rect 934 75216 940 75268
rect 992 75256 998 75268
rect 1964 75256 1992 75287
rect 2038 75284 2044 75336
rect 2096 75324 2102 75336
rect 2314 75324 2320 75336
rect 2096 75296 2141 75324
rect 2275 75296 2320 75324
rect 2096 75284 2102 75296
rect 2314 75284 2320 75296
rect 2372 75284 2378 75336
rect 2774 75324 2780 75336
rect 2735 75296 2780 75324
rect 2774 75284 2780 75296
rect 2832 75284 2838 75336
rect 9950 75324 9956 75336
rect 6886 75296 9956 75324
rect 992 75228 1992 75256
rect 992 75216 998 75228
rect 1964 75188 1992 75228
rect 2133 75259 2191 75265
rect 2133 75225 2145 75259
rect 2179 75256 2191 75259
rect 6886 75256 6914 75296
rect 9950 75284 9956 75296
rect 10008 75284 10014 75336
rect 10134 75324 10140 75336
rect 10095 75296 10140 75324
rect 10134 75284 10140 75296
rect 10192 75284 10198 75336
rect 2179 75228 6914 75256
rect 2179 75225 2191 75228
rect 2133 75219 2191 75225
rect 2590 75188 2596 75200
rect 1964 75160 2596 75188
rect 2590 75148 2596 75160
rect 2648 75148 2654 75200
rect 2961 75191 3019 75197
rect 2961 75157 2973 75191
rect 3007 75188 3019 75191
rect 4614 75188 4620 75200
rect 3007 75160 4620 75188
rect 3007 75157 3019 75160
rect 2961 75151 3019 75157
rect 4614 75148 4620 75160
rect 4672 75148 4678 75200
rect 9858 75148 9864 75200
rect 9916 75188 9922 75200
rect 9953 75191 10011 75197
rect 9953 75188 9965 75191
rect 9916 75160 9965 75188
rect 9916 75148 9922 75160
rect 9953 75157 9965 75160
rect 9999 75157 10011 75191
rect 9953 75151 10011 75157
rect 1104 75098 10856 75120
rect 1104 75046 4213 75098
rect 4265 75046 4277 75098
rect 4329 75046 4341 75098
rect 4393 75046 4405 75098
rect 4457 75046 4469 75098
rect 4521 75046 7477 75098
rect 7529 75046 7541 75098
rect 7593 75046 7605 75098
rect 7657 75046 7669 75098
rect 7721 75046 7733 75098
rect 7785 75046 10856 75098
rect 1104 75024 10856 75046
rect 9674 74984 9680 74996
rect 2148 74956 9680 74984
rect 934 74808 940 74860
rect 992 74848 998 74860
rect 2148 74857 2176 74956
rect 9674 74944 9680 74956
rect 9732 74944 9738 74996
rect 2866 74916 2872 74928
rect 2240 74888 2872 74916
rect 1897 74851 1955 74857
rect 1897 74848 1909 74851
rect 992 74820 1909 74848
rect 992 74808 998 74820
rect 1897 74817 1909 74820
rect 1943 74817 1955 74851
rect 1897 74811 1955 74817
rect 2041 74851 2099 74857
rect 2041 74817 2053 74851
rect 2087 74817 2099 74851
rect 2041 74811 2099 74817
rect 2133 74851 2191 74857
rect 2133 74817 2145 74851
rect 2179 74817 2191 74851
rect 2133 74811 2191 74817
rect 2056 74780 2084 74811
rect 2240 74780 2268 74888
rect 2866 74876 2872 74888
rect 2924 74876 2930 74928
rect 3142 74916 3148 74928
rect 3103 74888 3148 74916
rect 3142 74876 3148 74888
rect 3200 74876 3206 74928
rect 3237 74919 3295 74925
rect 3237 74885 3249 74919
rect 3283 74916 3295 74919
rect 5534 74916 5540 74928
rect 3283 74888 5540 74916
rect 3283 74885 3295 74888
rect 3237 74879 3295 74885
rect 5534 74876 5540 74888
rect 5592 74876 5598 74928
rect 2314 74808 2320 74860
rect 2372 74848 2378 74860
rect 2372 74820 2465 74848
rect 2372 74808 2378 74820
rect 2590 74808 2596 74860
rect 2648 74848 2654 74860
rect 3001 74851 3059 74857
rect 3001 74848 3013 74851
rect 2648 74820 3013 74848
rect 2648 74808 2654 74820
rect 3001 74817 3013 74820
rect 3047 74817 3059 74851
rect 3001 74811 3059 74817
rect 3421 74851 3479 74857
rect 3421 74817 3433 74851
rect 3467 74848 3479 74851
rect 5166 74848 5172 74860
rect 3467 74820 5172 74848
rect 3467 74817 3479 74820
rect 3421 74811 3479 74817
rect 2056 74752 2268 74780
rect 2332 74780 2360 74808
rect 3436 74780 3464 74811
rect 5166 74808 5172 74820
rect 5224 74808 5230 74860
rect 2332 74752 3464 74780
rect 1765 74715 1823 74721
rect 1765 74681 1777 74715
rect 1811 74712 1823 74715
rect 3694 74712 3700 74724
rect 1811 74684 3700 74712
rect 1811 74681 1823 74684
rect 1765 74675 1823 74681
rect 3694 74672 3700 74684
rect 3752 74672 3758 74724
rect 2869 74647 2927 74653
rect 2869 74613 2881 74647
rect 2915 74644 2927 74647
rect 2958 74644 2964 74656
rect 2915 74616 2964 74644
rect 2915 74613 2927 74616
rect 2869 74607 2927 74613
rect 2958 74604 2964 74616
rect 3016 74604 3022 74656
rect 1104 74554 10856 74576
rect 1104 74502 2582 74554
rect 2634 74502 2646 74554
rect 2698 74502 2710 74554
rect 2762 74502 2774 74554
rect 2826 74502 2838 74554
rect 2890 74502 5845 74554
rect 5897 74502 5909 74554
rect 5961 74502 5973 74554
rect 6025 74502 6037 74554
rect 6089 74502 6101 74554
rect 6153 74502 9109 74554
rect 9161 74502 9173 74554
rect 9225 74502 9237 74554
rect 9289 74502 9301 74554
rect 9353 74502 9365 74554
rect 9417 74502 10856 74554
rect 1104 74480 10856 74502
rect 2225 74375 2283 74381
rect 2225 74341 2237 74375
rect 2271 74372 2283 74375
rect 8294 74372 8300 74384
rect 2271 74344 8300 74372
rect 2271 74341 2283 74344
rect 2225 74335 2283 74341
rect 8294 74332 8300 74344
rect 8352 74332 8358 74384
rect 2590 74264 2596 74316
rect 2648 74304 2654 74316
rect 3510 74304 3516 74316
rect 2648 74276 3516 74304
rect 2648 74264 2654 74276
rect 3510 74264 3516 74276
rect 3568 74264 3574 74316
rect 1302 74196 1308 74248
rect 1360 74236 1366 74248
rect 1397 74239 1455 74245
rect 1397 74236 1409 74239
rect 1360 74208 1409 74236
rect 1360 74196 1366 74208
rect 1397 74205 1409 74208
rect 1443 74205 1455 74239
rect 1397 74199 1455 74205
rect 2314 74196 2320 74248
rect 2372 74245 2378 74248
rect 2372 74239 2415 74245
rect 2403 74205 2415 74239
rect 2372 74199 2415 74205
rect 2372 74196 2378 74199
rect 2498 74196 2504 74248
rect 2556 74236 2562 74248
rect 2774 74236 2780 74248
rect 2556 74208 2601 74236
rect 2735 74208 2780 74236
rect 2556 74196 2562 74208
rect 2774 74196 2780 74208
rect 2832 74196 2838 74248
rect 2866 74196 2872 74248
rect 2924 74236 2930 74248
rect 3973 74239 4031 74245
rect 3973 74236 3985 74239
rect 2924 74208 3985 74236
rect 2924 74196 2930 74208
rect 3973 74205 3985 74208
rect 4019 74205 4031 74239
rect 10134 74236 10140 74248
rect 10095 74208 10140 74236
rect 3973 74199 4031 74205
rect 10134 74196 10140 74208
rect 10192 74196 10198 74248
rect 2593 74171 2651 74177
rect 2593 74137 2605 74171
rect 2639 74168 2651 74171
rect 9766 74168 9772 74180
rect 2639 74140 9772 74168
rect 2639 74137 2651 74140
rect 2593 74131 2651 74137
rect 9766 74128 9772 74140
rect 9824 74128 9830 74180
rect 1581 74103 1639 74109
rect 1581 74069 1593 74103
rect 1627 74100 1639 74103
rect 1670 74100 1676 74112
rect 1627 74072 1676 74100
rect 1627 74069 1639 74072
rect 1581 74063 1639 74069
rect 1670 74060 1676 74072
rect 1728 74060 1734 74112
rect 3789 74103 3847 74109
rect 3789 74069 3801 74103
rect 3835 74100 3847 74103
rect 3970 74100 3976 74112
rect 3835 74072 3976 74100
rect 3835 74069 3847 74072
rect 3789 74063 3847 74069
rect 3970 74060 3976 74072
rect 4028 74060 4034 74112
rect 9950 74100 9956 74112
rect 9911 74072 9956 74100
rect 9950 74060 9956 74072
rect 10008 74060 10014 74112
rect 1104 74010 10856 74032
rect 1104 73958 4213 74010
rect 4265 73958 4277 74010
rect 4329 73958 4341 74010
rect 4393 73958 4405 74010
rect 4457 73958 4469 74010
rect 4521 73958 7477 74010
rect 7529 73958 7541 74010
rect 7593 73958 7605 74010
rect 7657 73958 7669 74010
rect 7721 73958 7733 74010
rect 7785 73958 10856 74010
rect 1104 73936 10856 73958
rect 2406 73856 2412 73908
rect 2464 73896 2470 73908
rect 2464 73868 2544 73896
rect 2464 73856 2470 73868
rect 2516 73837 2544 73868
rect 2501 73831 2559 73837
rect 2501 73797 2513 73831
rect 2547 73797 2559 73831
rect 2501 73791 2559 73797
rect 2593 73831 2651 73837
rect 2593 73797 2605 73831
rect 2639 73828 2651 73831
rect 9858 73828 9864 73840
rect 2639 73800 9864 73828
rect 2639 73797 2651 73800
rect 2593 73791 2651 73797
rect 9858 73788 9864 73800
rect 9916 73788 9922 73840
rect 1394 73760 1400 73772
rect 1355 73732 1400 73760
rect 1394 73720 1400 73732
rect 1452 73720 1458 73772
rect 2314 73720 2320 73772
rect 2372 73769 2378 73772
rect 2372 73763 2415 73769
rect 2403 73729 2415 73763
rect 2774 73760 2780 73772
rect 2687 73732 2780 73760
rect 2372 73723 2415 73729
rect 2372 73720 2378 73723
rect 2774 73720 2780 73732
rect 2832 73760 2838 73772
rect 3050 73760 3056 73772
rect 2832 73732 3056 73760
rect 2832 73720 2838 73732
rect 3050 73720 3056 73732
rect 3108 73720 3114 73772
rect 1581 73627 1639 73633
rect 1581 73593 1593 73627
rect 1627 73624 1639 73627
rect 2406 73624 2412 73636
rect 1627 73596 2412 73624
rect 1627 73593 1639 73596
rect 1581 73587 1639 73593
rect 2406 73584 2412 73596
rect 2464 73584 2470 73636
rect 2225 73559 2283 73565
rect 2225 73525 2237 73559
rect 2271 73556 2283 73559
rect 4982 73556 4988 73568
rect 2271 73528 4988 73556
rect 2271 73525 2283 73528
rect 2225 73519 2283 73525
rect 4982 73516 4988 73528
rect 5040 73516 5046 73568
rect 1104 73466 10856 73488
rect 1104 73414 2582 73466
rect 2634 73414 2646 73466
rect 2698 73414 2710 73466
rect 2762 73414 2774 73466
rect 2826 73414 2838 73466
rect 2890 73414 5845 73466
rect 5897 73414 5909 73466
rect 5961 73414 5973 73466
rect 6025 73414 6037 73466
rect 6089 73414 6101 73466
rect 6153 73414 9109 73466
rect 9161 73414 9173 73466
rect 9225 73414 9237 73466
rect 9289 73414 9301 73466
rect 9353 73414 9365 73466
rect 9417 73414 10856 73466
rect 1104 73392 10856 73414
rect 2225 73287 2283 73293
rect 2225 73253 2237 73287
rect 2271 73253 2283 73287
rect 2225 73247 2283 73253
rect 2240 73216 2268 73247
rect 2240 73188 3188 73216
rect 1302 73108 1308 73160
rect 1360 73148 1366 73160
rect 1397 73151 1455 73157
rect 1397 73148 1409 73151
rect 1360 73120 1409 73148
rect 1360 73108 1366 73120
rect 1397 73117 1409 73120
rect 1443 73117 1455 73151
rect 1397 73111 1455 73117
rect 2314 73108 2320 73160
rect 2372 73157 2378 73160
rect 2372 73151 2415 73157
rect 2403 73117 2415 73151
rect 2372 73111 2415 73117
rect 2777 73151 2835 73157
rect 2777 73117 2789 73151
rect 2823 73148 2835 73151
rect 3050 73148 3056 73160
rect 2823 73120 3056 73148
rect 2823 73117 2835 73120
rect 2777 73111 2835 73117
rect 2372 73108 2378 73111
rect 3050 73108 3056 73120
rect 3108 73108 3114 73160
rect 3160 73148 3188 73188
rect 5534 73148 5540 73160
rect 3160 73120 5540 73148
rect 5534 73108 5540 73120
rect 5592 73108 5598 73160
rect 9950 73148 9956 73160
rect 6886 73120 9956 73148
rect 2130 73040 2136 73092
rect 2188 73080 2194 73092
rect 2501 73083 2559 73089
rect 2501 73080 2513 73083
rect 2188 73052 2513 73080
rect 2188 73040 2194 73052
rect 2501 73049 2513 73052
rect 2547 73049 2559 73083
rect 2501 73043 2559 73049
rect 2593 73083 2651 73089
rect 2593 73049 2605 73083
rect 2639 73080 2651 73083
rect 6886 73080 6914 73120
rect 9950 73108 9956 73120
rect 10008 73108 10014 73160
rect 10134 73148 10140 73160
rect 10095 73120 10140 73148
rect 10134 73108 10140 73120
rect 10192 73108 10198 73160
rect 2639 73052 6914 73080
rect 2639 73049 2651 73052
rect 2593 73043 2651 73049
rect 1581 73015 1639 73021
rect 1581 72981 1593 73015
rect 1627 73012 1639 73015
rect 3142 73012 3148 73024
rect 1627 72984 3148 73012
rect 1627 72981 1639 72984
rect 1581 72975 1639 72981
rect 3142 72972 3148 72984
rect 3200 72972 3206 73024
rect 8386 72972 8392 73024
rect 8444 73012 8450 73024
rect 9953 73015 10011 73021
rect 9953 73012 9965 73015
rect 8444 72984 9965 73012
rect 8444 72972 8450 72984
rect 9953 72981 9965 72984
rect 9999 72981 10011 73015
rect 9953 72975 10011 72981
rect 1104 72922 10856 72944
rect 1104 72870 4213 72922
rect 4265 72870 4277 72922
rect 4329 72870 4341 72922
rect 4393 72870 4405 72922
rect 4457 72870 4469 72922
rect 4521 72870 7477 72922
rect 7529 72870 7541 72922
rect 7593 72870 7605 72922
rect 7657 72870 7669 72922
rect 7721 72870 7733 72922
rect 7785 72870 10856 72922
rect 1104 72848 10856 72870
rect 1854 72768 1860 72820
rect 1912 72808 1918 72820
rect 2130 72808 2136 72820
rect 1912 72780 2136 72808
rect 1912 72768 1918 72780
rect 2130 72768 2136 72780
rect 2188 72768 2194 72820
rect 1210 72632 1216 72684
rect 1268 72672 1274 72684
rect 1397 72675 1455 72681
rect 1397 72672 1409 72675
rect 1268 72644 1409 72672
rect 1268 72632 1274 72644
rect 1397 72641 1409 72644
rect 1443 72641 1455 72675
rect 2038 72672 2044 72684
rect 1999 72644 2044 72672
rect 1397 72635 1455 72641
rect 2038 72632 2044 72644
rect 2096 72632 2102 72684
rect 1581 72471 1639 72477
rect 1581 72437 1593 72471
rect 1627 72468 1639 72471
rect 1762 72468 1768 72480
rect 1627 72440 1768 72468
rect 1627 72437 1639 72440
rect 1581 72431 1639 72437
rect 1762 72428 1768 72440
rect 1820 72428 1826 72480
rect 1854 72428 1860 72480
rect 1912 72468 1918 72480
rect 2225 72471 2283 72477
rect 2225 72468 2237 72471
rect 1912 72440 2237 72468
rect 1912 72428 1918 72440
rect 2225 72437 2237 72440
rect 2271 72437 2283 72471
rect 2225 72431 2283 72437
rect 1104 72378 10856 72400
rect 1104 72326 2582 72378
rect 2634 72326 2646 72378
rect 2698 72326 2710 72378
rect 2762 72326 2774 72378
rect 2826 72326 2838 72378
rect 2890 72326 5845 72378
rect 5897 72326 5909 72378
rect 5961 72326 5973 72378
rect 6025 72326 6037 72378
rect 6089 72326 6101 72378
rect 6153 72326 9109 72378
rect 9161 72326 9173 72378
rect 9225 72326 9237 72378
rect 9289 72326 9301 72378
rect 9353 72326 9365 72378
rect 9417 72326 10856 72378
rect 1104 72304 10856 72326
rect 1026 72156 1032 72208
rect 1084 72196 1090 72208
rect 2225 72199 2283 72205
rect 2225 72196 2237 72199
rect 1084 72168 2237 72196
rect 1084 72156 1090 72168
rect 2225 72165 2237 72168
rect 2271 72165 2283 72199
rect 2225 72159 2283 72165
rect 1394 72060 1400 72072
rect 1355 72032 1400 72060
rect 1394 72020 1400 72032
rect 1452 72020 1458 72072
rect 1486 72020 1492 72072
rect 1544 72020 1550 72072
rect 2038 72020 2044 72072
rect 2096 72060 2102 72072
rect 2314 72060 2320 72072
rect 2372 72069 2378 72072
rect 2372 72063 2415 72069
rect 2096 72032 2320 72060
rect 2096 72020 2102 72032
rect 2314 72020 2320 72032
rect 2403 72029 2415 72063
rect 2372 72023 2415 72029
rect 2777 72063 2835 72069
rect 2777 72029 2789 72063
rect 2823 72060 2835 72063
rect 3050 72060 3056 72072
rect 2823 72032 3056 72060
rect 2823 72029 2835 72032
rect 2777 72023 2835 72029
rect 2372 72020 2378 72023
rect 3050 72020 3056 72032
rect 3108 72020 3114 72072
rect 10134 72060 10140 72072
rect 10095 72032 10140 72060
rect 10134 72020 10140 72032
rect 10192 72020 10198 72072
rect 1504 71992 1532 72020
rect 1504 71964 2176 71992
rect 1486 71884 1492 71936
rect 1544 71924 1550 71936
rect 1581 71927 1639 71933
rect 1581 71924 1593 71927
rect 1544 71896 1593 71924
rect 1544 71884 1550 71896
rect 1581 71893 1593 71896
rect 1627 71893 1639 71927
rect 2148 71924 2176 71964
rect 2222 71952 2228 72004
rect 2280 71992 2286 72004
rect 2501 71995 2559 72001
rect 2501 71992 2513 71995
rect 2280 71964 2513 71992
rect 2280 71952 2286 71964
rect 2501 71961 2513 71964
rect 2547 71961 2559 71995
rect 2501 71955 2559 71961
rect 2593 71995 2651 72001
rect 2593 71961 2605 71995
rect 2639 71992 2651 71995
rect 8386 71992 8392 72004
rect 2639 71964 8392 71992
rect 2639 71961 2651 71964
rect 2593 71955 2651 71961
rect 8386 71952 8392 71964
rect 8444 71952 8450 72004
rect 2314 71924 2320 71936
rect 2148 71896 2320 71924
rect 1581 71887 1639 71893
rect 2314 71884 2320 71896
rect 2372 71884 2378 71936
rect 9950 71924 9956 71936
rect 9911 71896 9956 71924
rect 9950 71884 9956 71896
rect 10008 71884 10014 71936
rect 1104 71834 10856 71856
rect 1104 71782 4213 71834
rect 4265 71782 4277 71834
rect 4329 71782 4341 71834
rect 4393 71782 4405 71834
rect 4457 71782 4469 71834
rect 4521 71782 7477 71834
rect 7529 71782 7541 71834
rect 7593 71782 7605 71834
rect 7657 71782 7669 71834
rect 7721 71782 7733 71834
rect 7785 71782 10856 71834
rect 1104 71760 10856 71782
rect 1578 71612 1584 71664
rect 1636 71652 1642 71664
rect 2501 71655 2559 71661
rect 2501 71652 2513 71655
rect 1636 71624 2513 71652
rect 1636 71612 1642 71624
rect 2501 71621 2513 71624
rect 2547 71621 2559 71655
rect 2501 71615 2559 71621
rect 2593 71655 2651 71661
rect 2593 71621 2605 71655
rect 2639 71652 2651 71655
rect 9950 71652 9956 71664
rect 2639 71624 9956 71652
rect 2639 71621 2651 71624
rect 2593 71615 2651 71621
rect 9950 71612 9956 71624
rect 10008 71612 10014 71664
rect 1302 71544 1308 71596
rect 1360 71584 1366 71596
rect 1397 71587 1455 71593
rect 1397 71584 1409 71587
rect 1360 71556 1409 71584
rect 1360 71544 1366 71556
rect 1397 71553 1409 71556
rect 1443 71553 1455 71587
rect 1397 71547 1455 71553
rect 2038 71544 2044 71596
rect 2096 71584 2102 71596
rect 2357 71587 2415 71593
rect 2357 71584 2369 71587
rect 2096 71556 2369 71584
rect 2096 71544 2102 71556
rect 2357 71553 2369 71556
rect 2403 71553 2415 71587
rect 2357 71547 2415 71553
rect 2777 71587 2835 71593
rect 2777 71553 2789 71587
rect 2823 71584 2835 71587
rect 3050 71584 3056 71596
rect 2823 71556 3056 71584
rect 2823 71553 2835 71556
rect 2777 71547 2835 71553
rect 3050 71544 3056 71556
rect 3108 71544 3114 71596
rect 1578 71380 1584 71392
rect 1539 71352 1584 71380
rect 1578 71340 1584 71352
rect 1636 71340 1642 71392
rect 2225 71383 2283 71389
rect 2225 71349 2237 71383
rect 2271 71380 2283 71383
rect 3234 71380 3240 71392
rect 2271 71352 3240 71380
rect 2271 71349 2283 71352
rect 2225 71343 2283 71349
rect 3234 71340 3240 71352
rect 3292 71340 3298 71392
rect 1104 71290 10856 71312
rect 1104 71238 2582 71290
rect 2634 71238 2646 71290
rect 2698 71238 2710 71290
rect 2762 71238 2774 71290
rect 2826 71238 2838 71290
rect 2890 71238 5845 71290
rect 5897 71238 5909 71290
rect 5961 71238 5973 71290
rect 6025 71238 6037 71290
rect 6089 71238 6101 71290
rect 6153 71238 9109 71290
rect 9161 71238 9173 71290
rect 9225 71238 9237 71290
rect 9289 71238 9301 71290
rect 9353 71238 9365 71290
rect 9417 71238 10856 71290
rect 1104 71216 10856 71238
rect 382 71068 388 71120
rect 440 71108 446 71120
rect 1949 71111 2007 71117
rect 1949 71108 1961 71111
rect 440 71080 1961 71108
rect 440 71068 446 71080
rect 1949 71077 1961 71080
rect 1995 71077 2007 71111
rect 1949 71071 2007 71077
rect 2314 71068 2320 71120
rect 2372 71108 2378 71120
rect 2590 71108 2596 71120
rect 2372 71080 2596 71108
rect 2372 71068 2378 71080
rect 2590 71068 2596 71080
rect 2648 71068 2654 71120
rect 1394 70972 1400 70984
rect 1355 70944 1400 70972
rect 1394 70932 1400 70944
rect 1452 70932 1458 70984
rect 1817 70975 1875 70981
rect 1817 70941 1829 70975
rect 1863 70972 1875 70975
rect 2314 70972 2320 70984
rect 1863 70944 2320 70972
rect 1863 70941 1875 70944
rect 1817 70935 1875 70941
rect 2314 70932 2320 70944
rect 2372 70932 2378 70984
rect 2685 70975 2743 70981
rect 2685 70941 2697 70975
rect 2731 70972 2743 70975
rect 2774 70972 2780 70984
rect 2731 70944 2780 70972
rect 2731 70941 2743 70944
rect 2685 70935 2743 70941
rect 2774 70932 2780 70944
rect 2832 70932 2838 70984
rect 10134 70972 10140 70984
rect 10095 70944 10140 70972
rect 10134 70932 10140 70944
rect 10192 70932 10198 70984
rect 1581 70907 1639 70913
rect 1581 70873 1593 70907
rect 1627 70873 1639 70907
rect 1581 70867 1639 70873
rect 1673 70907 1731 70913
rect 1673 70873 1685 70907
rect 1719 70904 1731 70907
rect 1946 70904 1952 70916
rect 1719 70876 1952 70904
rect 1719 70873 1731 70876
rect 1673 70867 1731 70873
rect 1596 70836 1624 70867
rect 1946 70864 1952 70876
rect 2004 70864 2010 70916
rect 9858 70904 9864 70916
rect 2148 70876 9864 70904
rect 2148 70836 2176 70876
rect 9858 70864 9864 70876
rect 9916 70864 9922 70916
rect 1596 70808 2176 70836
rect 2222 70796 2228 70848
rect 2280 70836 2286 70848
rect 2501 70839 2559 70845
rect 2501 70836 2513 70839
rect 2280 70808 2513 70836
rect 2280 70796 2286 70808
rect 2501 70805 2513 70808
rect 2547 70805 2559 70839
rect 9950 70836 9956 70848
rect 9911 70808 9956 70836
rect 2501 70799 2559 70805
rect 9950 70796 9956 70808
rect 10008 70796 10014 70848
rect 1104 70746 10856 70768
rect 1104 70694 4213 70746
rect 4265 70694 4277 70746
rect 4329 70694 4341 70746
rect 4393 70694 4405 70746
rect 4457 70694 4469 70746
rect 4521 70694 7477 70746
rect 7529 70694 7541 70746
rect 7593 70694 7605 70746
rect 7657 70694 7669 70746
rect 7721 70694 7733 70746
rect 7785 70694 10856 70746
rect 1104 70672 10856 70694
rect 1394 70524 1400 70576
rect 1452 70524 1458 70576
rect 2590 70524 2596 70576
rect 2648 70564 2654 70576
rect 2869 70567 2927 70573
rect 2648 70536 2820 70564
rect 2648 70524 2654 70536
rect 1412 70496 1440 70524
rect 2685 70499 2743 70505
rect 2685 70496 2697 70499
rect 1412 70468 2697 70496
rect 2685 70465 2697 70468
rect 2731 70465 2743 70499
rect 2792 70496 2820 70536
rect 2869 70533 2881 70567
rect 2915 70564 2927 70567
rect 9950 70564 9956 70576
rect 2915 70536 9956 70564
rect 2915 70533 2927 70536
rect 2869 70527 2927 70533
rect 9950 70524 9956 70536
rect 10008 70524 10014 70576
rect 2961 70499 3019 70505
rect 2961 70496 2973 70499
rect 2792 70468 2973 70496
rect 2685 70459 2743 70465
rect 2961 70465 2973 70468
rect 3007 70465 3019 70499
rect 2961 70459 3019 70465
rect 3058 70499 3116 70505
rect 3058 70465 3070 70499
rect 3104 70496 3116 70499
rect 3326 70496 3332 70508
rect 3104 70468 3332 70496
rect 3104 70465 3116 70468
rect 3058 70459 3116 70465
rect 1210 70388 1216 70440
rect 1268 70428 1274 70440
rect 1397 70431 1455 70437
rect 1397 70428 1409 70431
rect 1268 70400 1409 70428
rect 1268 70388 1274 70400
rect 1397 70397 1409 70400
rect 1443 70397 1455 70431
rect 1397 70391 1455 70397
rect 1673 70431 1731 70437
rect 1673 70397 1685 70431
rect 1719 70428 1731 70431
rect 1946 70428 1952 70440
rect 1719 70400 1952 70428
rect 1719 70397 1731 70400
rect 1673 70391 1731 70397
rect 1946 70388 1952 70400
rect 2004 70388 2010 70440
rect 2314 70388 2320 70440
rect 2372 70428 2378 70440
rect 3068 70428 3096 70459
rect 3326 70456 3332 70468
rect 3384 70456 3390 70508
rect 5258 70428 5264 70440
rect 2372 70400 3096 70428
rect 3252 70400 5264 70428
rect 2372 70388 2378 70400
rect 3252 70369 3280 70400
rect 5258 70388 5264 70400
rect 5316 70388 5322 70440
rect 3237 70363 3295 70369
rect 3237 70329 3249 70363
rect 3283 70360 3295 70363
rect 3283 70332 3317 70360
rect 3283 70329 3295 70332
rect 3237 70323 3295 70329
rect 1104 70202 10856 70224
rect 1104 70150 2582 70202
rect 2634 70150 2646 70202
rect 2698 70150 2710 70202
rect 2762 70150 2774 70202
rect 2826 70150 2838 70202
rect 2890 70150 5845 70202
rect 5897 70150 5909 70202
rect 5961 70150 5973 70202
rect 6025 70150 6037 70202
rect 6089 70150 6101 70202
rect 6153 70150 9109 70202
rect 9161 70150 9173 70202
rect 9225 70150 9237 70202
rect 9289 70150 9301 70202
rect 9353 70150 9365 70202
rect 9417 70150 10856 70202
rect 1104 70128 10856 70150
rect 9858 70048 9864 70100
rect 9916 70088 9922 70100
rect 9953 70091 10011 70097
rect 9953 70088 9965 70091
rect 9916 70060 9965 70088
rect 9916 70048 9922 70060
rect 9953 70057 9965 70060
rect 9999 70057 10011 70091
rect 9953 70051 10011 70057
rect 1394 69980 1400 70032
rect 1452 70020 1458 70032
rect 1578 70020 1584 70032
rect 1452 69992 1584 70020
rect 1452 69980 1458 69992
rect 1578 69980 1584 69992
rect 1636 69980 1642 70032
rect 842 69912 848 69964
rect 900 69952 906 69964
rect 1673 69955 1731 69961
rect 1673 69952 1685 69955
rect 900 69924 1685 69952
rect 900 69912 906 69924
rect 1673 69921 1685 69924
rect 1719 69921 1731 69955
rect 1673 69915 1731 69921
rect 1394 69884 1400 69896
rect 1355 69856 1400 69884
rect 1394 69844 1400 69856
rect 1452 69844 1458 69896
rect 2866 69884 2872 69896
rect 2827 69856 2872 69884
rect 2866 69844 2872 69856
rect 2924 69844 2930 69896
rect 10134 69884 10140 69896
rect 10095 69856 10140 69884
rect 10134 69844 10140 69856
rect 10192 69844 10198 69896
rect 2222 69708 2228 69760
rect 2280 69748 2286 69760
rect 2685 69751 2743 69757
rect 2685 69748 2697 69751
rect 2280 69720 2697 69748
rect 2280 69708 2286 69720
rect 2685 69717 2697 69720
rect 2731 69717 2743 69751
rect 2685 69711 2743 69717
rect 1104 69658 10856 69680
rect 1104 69606 4213 69658
rect 4265 69606 4277 69658
rect 4329 69606 4341 69658
rect 4393 69606 4405 69658
rect 4457 69606 4469 69658
rect 4521 69606 7477 69658
rect 7529 69606 7541 69658
rect 7593 69606 7605 69658
rect 7657 69606 7669 69658
rect 7721 69606 7733 69658
rect 7785 69606 10856 69658
rect 1104 69584 10856 69606
rect 2038 69436 2044 69488
rect 2096 69476 2102 69488
rect 2096 69448 2774 69476
rect 2096 69436 2102 69448
rect 2746 69408 2774 69448
rect 3050 69436 3056 69488
rect 3108 69476 3114 69488
rect 3108 69448 4476 69476
rect 3108 69436 3114 69448
rect 4448 69417 4476 69448
rect 3145 69411 3203 69417
rect 3145 69408 3157 69411
rect 2746 69380 3157 69408
rect 3145 69377 3157 69380
rect 3191 69377 3203 69411
rect 3145 69371 3203 69377
rect 4433 69411 4491 69417
rect 4433 69377 4445 69411
rect 4479 69377 4491 69411
rect 4433 69371 4491 69377
rect 1302 69300 1308 69352
rect 1360 69340 1366 69352
rect 1397 69343 1455 69349
rect 1397 69340 1409 69343
rect 1360 69312 1409 69340
rect 1360 69300 1366 69312
rect 1397 69309 1409 69312
rect 1443 69309 1455 69343
rect 1397 69303 1455 69309
rect 1673 69343 1731 69349
rect 1673 69309 1685 69343
rect 1719 69340 1731 69343
rect 2038 69340 2044 69352
rect 1719 69312 2044 69340
rect 1719 69309 1731 69312
rect 1673 69303 1731 69309
rect 2038 69300 2044 69312
rect 2096 69300 2102 69352
rect 2869 69343 2927 69349
rect 2869 69309 2881 69343
rect 2915 69340 2927 69343
rect 3050 69340 3056 69352
rect 2915 69312 3056 69340
rect 2915 69309 2927 69312
rect 2869 69303 2927 69309
rect 3050 69300 3056 69312
rect 3108 69300 3114 69352
rect 3418 69300 3424 69352
rect 3476 69340 3482 69352
rect 4157 69343 4215 69349
rect 4157 69340 4169 69343
rect 3476 69312 4169 69340
rect 3476 69300 3482 69312
rect 4157 69309 4169 69312
rect 4203 69309 4215 69343
rect 4157 69303 4215 69309
rect 1104 69114 10856 69136
rect 1104 69062 2582 69114
rect 2634 69062 2646 69114
rect 2698 69062 2710 69114
rect 2762 69062 2774 69114
rect 2826 69062 2838 69114
rect 2890 69062 5845 69114
rect 5897 69062 5909 69114
rect 5961 69062 5973 69114
rect 6025 69062 6037 69114
rect 6089 69062 6101 69114
rect 6153 69062 9109 69114
rect 9161 69062 9173 69114
rect 9225 69062 9237 69114
rect 9289 69062 9301 69114
rect 9353 69062 9365 69114
rect 9417 69062 10856 69114
rect 1104 69040 10856 69062
rect 1578 68892 1584 68944
rect 1636 68932 1642 68944
rect 2314 68932 2320 68944
rect 1636 68904 2320 68932
rect 1636 68892 1642 68904
rect 2314 68892 2320 68904
rect 2372 68932 2378 68944
rect 3878 68932 3884 68944
rect 2372 68904 2774 68932
rect 3839 68904 3884 68932
rect 2372 68892 2378 68904
rect 2746 68864 2774 68904
rect 3878 68892 3884 68904
rect 3936 68892 3942 68944
rect 2746 68836 4476 68864
rect 1394 68796 1400 68808
rect 1355 68768 1400 68796
rect 1394 68756 1400 68768
rect 1452 68756 1458 68808
rect 1578 68756 1584 68808
rect 1636 68796 1642 68808
rect 1673 68799 1731 68805
rect 1673 68796 1685 68799
rect 1636 68768 1685 68796
rect 1636 68756 1642 68768
rect 1673 68765 1685 68768
rect 1719 68765 1731 68799
rect 1673 68759 1731 68765
rect 3326 68756 3332 68808
rect 3384 68796 3390 68808
rect 4448 68805 4476 68836
rect 4013 68799 4071 68805
rect 4013 68796 4025 68799
rect 3384 68768 4025 68796
rect 3384 68756 3390 68768
rect 4013 68765 4025 68768
rect 4059 68765 4071 68799
rect 4013 68759 4071 68765
rect 4433 68799 4491 68805
rect 4433 68765 4445 68799
rect 4479 68796 4491 68799
rect 4706 68796 4712 68808
rect 4479 68768 4712 68796
rect 4479 68765 4491 68768
rect 4433 68759 4491 68765
rect 4706 68756 4712 68768
rect 4764 68756 4770 68808
rect 10134 68796 10140 68808
rect 10095 68768 10140 68796
rect 10134 68756 10140 68768
rect 10192 68756 10198 68808
rect 2498 68688 2504 68740
rect 2556 68728 2562 68740
rect 4157 68731 4215 68737
rect 4157 68728 4169 68731
rect 2556 68700 4169 68728
rect 2556 68688 2562 68700
rect 4157 68697 4169 68700
rect 4203 68697 4215 68731
rect 4157 68691 4215 68697
rect 4249 68731 4307 68737
rect 4249 68697 4261 68731
rect 4295 68728 4307 68731
rect 4295 68700 9996 68728
rect 4295 68697 4307 68700
rect 4249 68691 4307 68697
rect 1762 68620 1768 68672
rect 1820 68660 1826 68672
rect 2590 68660 2596 68672
rect 1820 68632 2596 68660
rect 1820 68620 1826 68632
rect 2590 68620 2596 68632
rect 2648 68620 2654 68672
rect 9968 68669 9996 68700
rect 9953 68663 10011 68669
rect 9953 68629 9965 68663
rect 9999 68629 10011 68663
rect 9953 68623 10011 68629
rect 1104 68570 10856 68592
rect 1104 68518 4213 68570
rect 4265 68518 4277 68570
rect 4329 68518 4341 68570
rect 4393 68518 4405 68570
rect 4457 68518 4469 68570
rect 4521 68518 7477 68570
rect 7529 68518 7541 68570
rect 7593 68518 7605 68570
rect 7657 68518 7669 68570
rect 7721 68518 7733 68570
rect 7785 68518 10856 68570
rect 1104 68496 10856 68518
rect 1854 68416 1860 68468
rect 1912 68456 1918 68468
rect 2222 68456 2228 68468
rect 1912 68428 2228 68456
rect 1912 68416 1918 68428
rect 2222 68416 2228 68428
rect 2280 68416 2286 68468
rect 3050 68388 3056 68400
rect 1688 68360 2452 68388
rect 1688 68329 1716 68360
rect 1668 68323 1726 68329
rect 1668 68289 1680 68323
rect 1714 68289 1726 68323
rect 1668 68283 1726 68289
rect 1764 68323 1822 68329
rect 1764 68289 1776 68323
rect 1810 68289 1822 68323
rect 1764 68283 1822 68289
rect 1857 68323 1915 68329
rect 1857 68289 1869 68323
rect 1903 68320 1915 68323
rect 2041 68323 2099 68329
rect 1903 68292 1992 68320
rect 1903 68289 1915 68292
rect 1857 68283 1915 68289
rect 1486 68212 1492 68264
rect 1544 68212 1550 68264
rect 1780 68252 1808 68283
rect 1780 68224 1900 68252
rect 1504 68184 1532 68212
rect 1504 68156 1808 68184
rect 1780 68128 1808 68156
rect 1486 68116 1492 68128
rect 1447 68088 1492 68116
rect 1486 68076 1492 68088
rect 1544 68076 1550 68128
rect 1762 68076 1768 68128
rect 1820 68076 1826 68128
rect 1872 68116 1900 68224
rect 1964 68184 1992 68292
rect 2041 68289 2053 68323
rect 2087 68320 2099 68323
rect 2314 68320 2320 68332
rect 2087 68292 2320 68320
rect 2087 68289 2099 68292
rect 2041 68283 2099 68289
rect 2314 68280 2320 68292
rect 2372 68280 2378 68332
rect 2424 68252 2452 68360
rect 2746 68360 3056 68388
rect 2593 68323 2651 68329
rect 2593 68289 2605 68323
rect 2639 68320 2651 68323
rect 2746 68320 2774 68360
rect 3050 68348 3056 68360
rect 3108 68388 3114 68400
rect 3510 68388 3516 68400
rect 3108 68360 3516 68388
rect 3108 68348 3114 68360
rect 3510 68348 3516 68360
rect 3568 68348 3574 68400
rect 4249 68391 4307 68397
rect 4249 68357 4261 68391
rect 4295 68388 4307 68391
rect 4614 68388 4620 68400
rect 4295 68360 4620 68388
rect 4295 68357 4307 68360
rect 4249 68351 4307 68357
rect 4614 68348 4620 68360
rect 4672 68348 4678 68400
rect 2639 68292 2774 68320
rect 2869 68323 2927 68329
rect 2639 68289 2651 68292
rect 2593 68283 2651 68289
rect 2869 68289 2881 68323
rect 2915 68320 2927 68323
rect 3326 68320 3332 68332
rect 2915 68292 3332 68320
rect 2915 68289 2927 68292
rect 2869 68283 2927 68289
rect 2884 68252 2912 68283
rect 3326 68280 3332 68292
rect 3384 68320 3390 68332
rect 4105 68323 4163 68329
rect 4105 68320 4117 68323
rect 3384 68292 4117 68320
rect 3384 68280 3390 68292
rect 4105 68289 4117 68292
rect 4151 68289 4163 68323
rect 4105 68283 4163 68289
rect 4338 68280 4344 68332
rect 4396 68320 4402 68332
rect 4525 68323 4583 68329
rect 4396 68292 4441 68320
rect 4396 68280 4402 68292
rect 4525 68289 4537 68323
rect 4571 68320 4583 68323
rect 4706 68320 4712 68332
rect 4571 68292 4712 68320
rect 4571 68289 4583 68292
rect 4525 68283 4583 68289
rect 4706 68280 4712 68292
rect 4764 68280 4770 68332
rect 2424 68224 2912 68252
rect 9950 68184 9956 68196
rect 1964 68156 9956 68184
rect 9950 68144 9956 68156
rect 10008 68144 10014 68196
rect 2130 68116 2136 68128
rect 1872 68088 2136 68116
rect 2130 68076 2136 68088
rect 2188 68076 2194 68128
rect 3973 68119 4031 68125
rect 3973 68085 3985 68119
rect 4019 68116 4031 68119
rect 8386 68116 8392 68128
rect 4019 68088 8392 68116
rect 4019 68085 4031 68088
rect 3973 68079 4031 68085
rect 8386 68076 8392 68088
rect 8444 68076 8450 68128
rect 1104 68026 10856 68048
rect 1104 67974 2582 68026
rect 2634 67974 2646 68026
rect 2698 67974 2710 68026
rect 2762 67974 2774 68026
rect 2826 67974 2838 68026
rect 2890 67974 5845 68026
rect 5897 67974 5909 68026
rect 5961 67974 5973 68026
rect 6025 67974 6037 68026
rect 6089 67974 6101 68026
rect 6153 67974 9109 68026
rect 9161 67974 9173 68026
rect 9225 67974 9237 68026
rect 9289 67974 9301 68026
rect 9353 67974 9365 68026
rect 9417 67974 10856 68026
rect 1104 67952 10856 67974
rect 1486 67872 1492 67924
rect 1544 67912 1550 67924
rect 1544 67884 2774 67912
rect 1544 67872 1550 67884
rect 2746 67844 2774 67884
rect 4338 67872 4344 67924
rect 4396 67912 4402 67924
rect 9953 67915 10011 67921
rect 9953 67912 9965 67915
rect 4396 67884 9965 67912
rect 4396 67872 4402 67884
rect 9953 67881 9965 67884
rect 9999 67881 10011 67915
rect 9953 67875 10011 67881
rect 6914 67844 6920 67856
rect 2746 67816 6920 67844
rect 6914 67804 6920 67816
rect 6972 67804 6978 67856
rect 2314 67736 2320 67788
rect 2372 67776 2378 67788
rect 2869 67779 2927 67785
rect 2869 67776 2881 67779
rect 2372 67748 2881 67776
rect 2372 67736 2378 67748
rect 2869 67745 2881 67748
rect 2915 67745 2927 67779
rect 2869 67739 2927 67745
rect 3145 67779 3203 67785
rect 3145 67745 3157 67779
rect 3191 67776 3203 67779
rect 3418 67776 3424 67788
rect 3191 67748 3424 67776
rect 3191 67745 3203 67748
rect 3145 67739 3203 67745
rect 3418 67736 3424 67748
rect 3476 67776 3482 67788
rect 3602 67776 3608 67788
rect 3476 67748 3608 67776
rect 3476 67736 3482 67748
rect 3602 67736 3608 67748
rect 3660 67736 3666 67788
rect 10137 67711 10195 67717
rect 10137 67677 10149 67711
rect 10183 67677 10195 67711
rect 10137 67671 10195 67677
rect 1670 67640 1676 67652
rect 1631 67612 1676 67640
rect 1670 67600 1676 67612
rect 1728 67600 1734 67652
rect 1857 67643 1915 67649
rect 1857 67609 1869 67643
rect 1903 67640 1915 67643
rect 4706 67640 4712 67652
rect 1903 67612 4712 67640
rect 1903 67609 1915 67612
rect 1857 67603 1915 67609
rect 4706 67600 4712 67612
rect 4764 67600 4770 67652
rect 10152 67584 10180 67671
rect 10134 67532 10140 67584
rect 10192 67532 10198 67584
rect 1104 67482 10856 67504
rect 1104 67430 4213 67482
rect 4265 67430 4277 67482
rect 4329 67430 4341 67482
rect 4393 67430 4405 67482
rect 4457 67430 4469 67482
rect 4521 67430 7477 67482
rect 7529 67430 7541 67482
rect 7593 67430 7605 67482
rect 7657 67430 7669 67482
rect 7721 67430 7733 67482
rect 7785 67430 10856 67482
rect 1104 67408 10856 67430
rect 1394 67232 1400 67244
rect 1355 67204 1400 67232
rect 1394 67192 1400 67204
rect 1452 67192 1458 67244
rect 1673 67167 1731 67173
rect 1673 67133 1685 67167
rect 1719 67133 1731 67167
rect 1673 67127 1731 67133
rect 1688 67040 1716 67127
rect 1670 66988 1676 67040
rect 1728 66988 1734 67040
rect 1104 66938 10856 66960
rect 1104 66886 2582 66938
rect 2634 66886 2646 66938
rect 2698 66886 2710 66938
rect 2762 66886 2774 66938
rect 2826 66886 2838 66938
rect 2890 66886 5845 66938
rect 5897 66886 5909 66938
rect 5961 66886 5973 66938
rect 6025 66886 6037 66938
rect 6089 66886 6101 66938
rect 6153 66886 9109 66938
rect 9161 66886 9173 66938
rect 9225 66886 9237 66938
rect 9289 66886 9301 66938
rect 9353 66886 9365 66938
rect 9417 66886 10856 66938
rect 1104 66864 10856 66886
rect 1394 66512 1400 66564
rect 1452 66552 1458 66564
rect 1949 66555 2007 66561
rect 1949 66552 1961 66555
rect 1452 66524 1961 66552
rect 1452 66512 1458 66524
rect 1949 66521 1961 66524
rect 1995 66521 2007 66555
rect 1949 66515 2007 66521
rect 2685 66555 2743 66561
rect 2685 66521 2697 66555
rect 2731 66552 2743 66555
rect 2774 66552 2780 66564
rect 2731 66524 2780 66552
rect 2731 66521 2743 66524
rect 2685 66515 2743 66521
rect 2774 66512 2780 66524
rect 2832 66512 2838 66564
rect 658 66444 664 66496
rect 716 66484 722 66496
rect 1857 66487 1915 66493
rect 1857 66484 1869 66487
rect 716 66456 1869 66484
rect 716 66444 722 66456
rect 1857 66453 1869 66456
rect 1903 66453 1915 66487
rect 1857 66447 1915 66453
rect 2593 66487 2651 66493
rect 2593 66453 2605 66487
rect 2639 66484 2651 66487
rect 3418 66484 3424 66496
rect 2639 66456 3424 66484
rect 2639 66453 2651 66456
rect 2593 66447 2651 66453
rect 3418 66444 3424 66456
rect 3476 66444 3482 66496
rect 1104 66394 10856 66416
rect 1104 66342 4213 66394
rect 4265 66342 4277 66394
rect 4329 66342 4341 66394
rect 4393 66342 4405 66394
rect 4457 66342 4469 66394
rect 4521 66342 7477 66394
rect 7529 66342 7541 66394
rect 7593 66342 7605 66394
rect 7657 66342 7669 66394
rect 7721 66342 7733 66394
rect 7785 66342 10856 66394
rect 1104 66320 10856 66342
rect 1946 66240 1952 66292
rect 2004 66280 2010 66292
rect 2130 66280 2136 66292
rect 2004 66252 2136 66280
rect 2004 66240 2010 66252
rect 2130 66240 2136 66252
rect 2188 66240 2194 66292
rect 9950 66280 9956 66292
rect 9911 66252 9956 66280
rect 9950 66240 9956 66252
rect 10008 66240 10014 66292
rect 1946 66144 1952 66156
rect 1907 66116 1952 66144
rect 1946 66104 1952 66116
rect 2004 66104 2010 66156
rect 2869 66147 2927 66153
rect 2869 66113 2881 66147
rect 2915 66144 2927 66147
rect 4062 66144 4068 66156
rect 2915 66116 4068 66144
rect 2915 66113 2927 66116
rect 2869 66107 2927 66113
rect 4062 66104 4068 66116
rect 4120 66104 4126 66156
rect 10134 66144 10140 66156
rect 10095 66116 10140 66144
rect 10134 66104 10140 66116
rect 10192 66104 10198 66156
rect 1765 66011 1823 66017
rect 1765 65977 1777 66011
rect 1811 66008 1823 66011
rect 8478 66008 8484 66020
rect 1811 65980 8484 66008
rect 1811 65977 1823 65980
rect 1765 65971 1823 65977
rect 8478 65968 8484 65980
rect 8536 65968 8542 66020
rect 3053 65943 3111 65949
rect 3053 65909 3065 65943
rect 3099 65940 3111 65943
rect 3142 65940 3148 65952
rect 3099 65912 3148 65940
rect 3099 65909 3111 65912
rect 3053 65903 3111 65909
rect 3142 65900 3148 65912
rect 3200 65900 3206 65952
rect 1104 65850 10856 65872
rect 1104 65798 2582 65850
rect 2634 65798 2646 65850
rect 2698 65798 2710 65850
rect 2762 65798 2774 65850
rect 2826 65798 2838 65850
rect 2890 65798 5845 65850
rect 5897 65798 5909 65850
rect 5961 65798 5973 65850
rect 6025 65798 6037 65850
rect 6089 65798 6101 65850
rect 6153 65798 9109 65850
rect 9161 65798 9173 65850
rect 9225 65798 9237 65850
rect 9289 65798 9301 65850
rect 9353 65798 9365 65850
rect 9417 65798 10856 65850
rect 1104 65776 10856 65798
rect 2314 65628 2320 65680
rect 2372 65668 2378 65680
rect 3050 65668 3056 65680
rect 2372 65640 3056 65668
rect 2372 65628 2378 65640
rect 3050 65628 3056 65640
rect 3108 65628 3114 65680
rect 2777 65535 2835 65541
rect 2777 65501 2789 65535
rect 2823 65532 2835 65535
rect 3786 65532 3792 65544
rect 2823 65504 3792 65532
rect 2823 65501 2835 65504
rect 2777 65495 2835 65501
rect 3786 65492 3792 65504
rect 3844 65492 3850 65544
rect 750 65424 756 65476
rect 808 65464 814 65476
rect 1765 65467 1823 65473
rect 1765 65464 1777 65467
rect 808 65436 1777 65464
rect 808 65424 814 65436
rect 1765 65433 1777 65436
rect 1811 65433 1823 65467
rect 1946 65464 1952 65476
rect 1907 65436 1952 65464
rect 1765 65427 1823 65433
rect 1946 65424 1952 65436
rect 2004 65424 2010 65476
rect 2593 65399 2651 65405
rect 2593 65365 2605 65399
rect 2639 65396 2651 65399
rect 3050 65396 3056 65408
rect 2639 65368 3056 65396
rect 2639 65365 2651 65368
rect 2593 65359 2651 65365
rect 3050 65356 3056 65368
rect 3108 65356 3114 65408
rect 1104 65306 10856 65328
rect 1104 65254 4213 65306
rect 4265 65254 4277 65306
rect 4329 65254 4341 65306
rect 4393 65254 4405 65306
rect 4457 65254 4469 65306
rect 4521 65254 7477 65306
rect 7529 65254 7541 65306
rect 7593 65254 7605 65306
rect 7657 65254 7669 65306
rect 7721 65254 7733 65306
rect 7785 65254 10856 65306
rect 1104 65232 10856 65254
rect 5074 65124 5080 65136
rect 1688 65096 5080 65124
rect 1688 65065 1716 65096
rect 5074 65084 5080 65096
rect 5132 65084 5138 65136
rect 1673 65059 1731 65065
rect 1673 65025 1685 65059
rect 1719 65025 1731 65059
rect 1673 65019 1731 65025
rect 1946 65016 1952 65068
rect 2004 65056 2010 65068
rect 2314 65056 2320 65068
rect 2004 65028 2320 65056
rect 2004 65016 2010 65028
rect 2314 65016 2320 65028
rect 2372 65016 2378 65068
rect 2777 65059 2835 65065
rect 2777 65025 2789 65059
rect 2823 65056 2835 65059
rect 3510 65056 3516 65068
rect 2823 65028 3516 65056
rect 2823 65025 2835 65028
rect 2777 65019 2835 65025
rect 3510 65016 3516 65028
rect 3568 65016 3574 65068
rect 10134 65056 10140 65068
rect 10095 65028 10140 65056
rect 10134 65016 10140 65028
rect 10192 65016 10198 65068
rect 1486 64920 1492 64932
rect 1447 64892 1492 64920
rect 1486 64880 1492 64892
rect 1544 64880 1550 64932
rect 934 64812 940 64864
rect 992 64852 998 64864
rect 2314 64852 2320 64864
rect 992 64824 2320 64852
rect 992 64812 998 64824
rect 2314 64812 2320 64824
rect 2372 64852 2378 64864
rect 2961 64855 3019 64861
rect 2961 64852 2973 64855
rect 2372 64824 2973 64852
rect 2372 64812 2378 64824
rect 2961 64821 2973 64824
rect 3007 64821 3019 64855
rect 9950 64852 9956 64864
rect 9911 64824 9956 64852
rect 2961 64815 3019 64821
rect 9950 64812 9956 64824
rect 10008 64812 10014 64864
rect 1104 64762 10856 64784
rect 1104 64710 2582 64762
rect 2634 64710 2646 64762
rect 2698 64710 2710 64762
rect 2762 64710 2774 64762
rect 2826 64710 2838 64762
rect 2890 64710 5845 64762
rect 5897 64710 5909 64762
rect 5961 64710 5973 64762
rect 6025 64710 6037 64762
rect 6089 64710 6101 64762
rect 6153 64710 9109 64762
rect 9161 64710 9173 64762
rect 9225 64710 9237 64762
rect 9289 64710 9301 64762
rect 9353 64710 9365 64762
rect 9417 64710 10856 64762
rect 1104 64688 10856 64710
rect 14 64540 20 64592
rect 72 64580 78 64592
rect 2133 64583 2191 64589
rect 2133 64580 2145 64583
rect 72 64552 2145 64580
rect 72 64540 78 64552
rect 2133 64549 2145 64552
rect 2179 64549 2191 64583
rect 2133 64543 2191 64549
rect 3970 64512 3976 64524
rect 2424 64484 3976 64512
rect 2314 64453 2320 64456
rect 2312 64444 2320 64453
rect 2275 64416 2320 64444
rect 2312 64407 2320 64416
rect 2314 64404 2320 64407
rect 2372 64404 2378 64456
rect 2424 64453 2452 64484
rect 3970 64472 3976 64484
rect 4028 64472 4034 64524
rect 2409 64447 2467 64453
rect 2409 64413 2421 64447
rect 2455 64413 2467 64447
rect 2409 64407 2467 64413
rect 2685 64447 2743 64453
rect 2685 64413 2697 64447
rect 2731 64444 2743 64447
rect 2774 64444 2780 64456
rect 2731 64416 2780 64444
rect 2731 64413 2743 64416
rect 2685 64407 2743 64413
rect 2774 64404 2780 64416
rect 2832 64404 2838 64456
rect 3326 64404 3332 64456
rect 3384 64444 3390 64456
rect 3789 64447 3847 64453
rect 3789 64444 3801 64447
rect 3384 64416 3801 64444
rect 3384 64404 3390 64416
rect 3789 64413 3801 64416
rect 3835 64413 3847 64447
rect 3789 64407 3847 64413
rect 2501 64379 2559 64385
rect 2501 64345 2513 64379
rect 2547 64376 2559 64379
rect 9950 64376 9956 64388
rect 2547 64348 9956 64376
rect 2547 64345 2559 64348
rect 2501 64339 2559 64345
rect 9950 64336 9956 64348
rect 10008 64336 10014 64388
rect 3970 64308 3976 64320
rect 3931 64280 3976 64308
rect 3970 64268 3976 64280
rect 4028 64268 4034 64320
rect 1104 64218 10856 64240
rect 1104 64166 4213 64218
rect 4265 64166 4277 64218
rect 4329 64166 4341 64218
rect 4393 64166 4405 64218
rect 4457 64166 4469 64218
rect 4521 64166 7477 64218
rect 7529 64166 7541 64218
rect 7593 64166 7605 64218
rect 7657 64166 7669 64218
rect 7721 64166 7733 64218
rect 7785 64166 10856 64218
rect 1104 64144 10856 64166
rect 9953 64107 10011 64113
rect 9953 64104 9965 64107
rect 2746 64076 9965 64104
rect 1394 63996 1400 64048
rect 1452 64036 1458 64048
rect 2501 64039 2559 64045
rect 2501 64036 2513 64039
rect 1452 64008 2513 64036
rect 1452 63996 1458 64008
rect 2501 64005 2513 64008
rect 2547 64005 2559 64039
rect 2501 63999 2559 64005
rect 2593 64039 2651 64045
rect 2593 64005 2605 64039
rect 2639 64036 2651 64039
rect 2746 64036 2774 64076
rect 9953 64073 9965 64076
rect 9999 64073 10011 64107
rect 9953 64067 10011 64073
rect 2639 64008 2774 64036
rect 2639 64005 2651 64008
rect 2593 63999 2651 64005
rect 934 63928 940 63980
rect 992 63968 998 63980
rect 1673 63971 1731 63977
rect 1673 63968 1685 63971
rect 992 63940 1685 63968
rect 992 63928 998 63940
rect 1673 63937 1685 63940
rect 1719 63937 1731 63971
rect 1673 63931 1731 63937
rect 2314 63928 2320 63980
rect 2372 63977 2378 63980
rect 2372 63971 2415 63977
rect 2403 63937 2415 63971
rect 2372 63931 2415 63937
rect 2372 63928 2378 63931
rect 2774 63928 2780 63980
rect 2832 63968 2838 63980
rect 3050 63968 3056 63980
rect 2832 63940 3056 63968
rect 2832 63928 2838 63940
rect 3050 63928 3056 63940
rect 3108 63928 3114 63980
rect 10134 63968 10140 63980
rect 10095 63940 10140 63968
rect 10134 63928 10140 63940
rect 10192 63928 10198 63980
rect 1394 63724 1400 63776
rect 1452 63764 1458 63776
rect 1489 63767 1547 63773
rect 1489 63764 1501 63767
rect 1452 63736 1501 63764
rect 1452 63724 1458 63736
rect 1489 63733 1501 63736
rect 1535 63733 1547 63767
rect 1489 63727 1547 63733
rect 2225 63767 2283 63773
rect 2225 63733 2237 63767
rect 2271 63764 2283 63767
rect 6730 63764 6736 63776
rect 2271 63736 6736 63764
rect 2271 63733 2283 63736
rect 2225 63727 2283 63733
rect 6730 63724 6736 63736
rect 6788 63724 6794 63776
rect 1104 63674 10856 63696
rect 1104 63622 2582 63674
rect 2634 63622 2646 63674
rect 2698 63622 2710 63674
rect 2762 63622 2774 63674
rect 2826 63622 2838 63674
rect 2890 63622 5845 63674
rect 5897 63622 5909 63674
rect 5961 63622 5973 63674
rect 6025 63622 6037 63674
rect 6089 63622 6101 63674
rect 6153 63622 9109 63674
rect 9161 63622 9173 63674
rect 9225 63622 9237 63674
rect 9289 63622 9301 63674
rect 9353 63622 9365 63674
rect 9417 63622 10856 63674
rect 1104 63600 10856 63622
rect 2409 63427 2467 63433
rect 2409 63393 2421 63427
rect 2455 63424 2467 63427
rect 3510 63424 3516 63436
rect 2455 63396 3516 63424
rect 2455 63393 2467 63396
rect 2409 63387 2467 63393
rect 3510 63384 3516 63396
rect 3568 63384 3574 63436
rect 1673 63359 1731 63365
rect 1673 63325 1685 63359
rect 1719 63325 1731 63359
rect 1673 63319 1731 63325
rect 3789 63359 3847 63365
rect 3789 63325 3801 63359
rect 3835 63356 3847 63359
rect 5718 63356 5724 63368
rect 3835 63328 5724 63356
rect 3835 63325 3847 63328
rect 3789 63319 3847 63325
rect 1688 63288 1716 63319
rect 5718 63316 5724 63328
rect 5776 63316 5782 63368
rect 7374 63288 7380 63300
rect 1688 63260 7380 63288
rect 7374 63248 7380 63260
rect 7432 63248 7438 63300
rect 1486 63220 1492 63232
rect 1447 63192 1492 63220
rect 1486 63180 1492 63192
rect 1544 63180 1550 63232
rect 2314 63180 2320 63232
rect 2372 63220 2378 63232
rect 2639 63223 2697 63229
rect 2639 63220 2651 63223
rect 2372 63192 2651 63220
rect 2372 63180 2378 63192
rect 2639 63189 2651 63192
rect 2685 63189 2697 63223
rect 3970 63220 3976 63232
rect 3931 63192 3976 63220
rect 2639 63183 2697 63189
rect 3970 63180 3976 63192
rect 4028 63180 4034 63232
rect 1104 63130 10856 63152
rect 1104 63078 4213 63130
rect 4265 63078 4277 63130
rect 4329 63078 4341 63130
rect 4393 63078 4405 63130
rect 4457 63078 4469 63130
rect 4521 63078 7477 63130
rect 7529 63078 7541 63130
rect 7593 63078 7605 63130
rect 7657 63078 7669 63130
rect 7721 63078 7733 63130
rect 7785 63078 10856 63130
rect 1104 63056 10856 63078
rect 2406 63016 2412 63028
rect 1964 62988 2412 63016
rect 1964 62957 1992 62988
rect 2406 62976 2412 62988
rect 2464 62976 2470 63028
rect 9953 63019 10011 63025
rect 9953 63016 9965 63019
rect 2746 62988 9965 63016
rect 1949 62951 2007 62957
rect 1949 62917 1961 62951
rect 1995 62917 2007 62951
rect 1949 62911 2007 62917
rect 2041 62951 2099 62957
rect 2041 62917 2053 62951
rect 2087 62948 2099 62951
rect 2746 62948 2774 62988
rect 9953 62985 9965 62988
rect 9999 62985 10011 63019
rect 9953 62979 10011 62985
rect 2087 62920 2774 62948
rect 2087 62917 2099 62920
rect 2041 62911 2099 62917
rect 1852 62883 1910 62889
rect 1852 62849 1864 62883
rect 1898 62880 1910 62883
rect 2225 62883 2283 62889
rect 1898 62852 2176 62880
rect 1898 62849 1910 62852
rect 1852 62843 1910 62849
rect 2148 62812 2176 62852
rect 2225 62849 2237 62883
rect 2271 62880 2283 62883
rect 2961 62883 3019 62889
rect 2961 62880 2973 62883
rect 2271 62852 2973 62880
rect 2271 62849 2283 62852
rect 2225 62843 2283 62849
rect 2961 62849 2973 62852
rect 3007 62880 3019 62883
rect 3050 62880 3056 62892
rect 3007 62852 3056 62880
rect 3007 62849 3019 62852
rect 2961 62843 3019 62849
rect 3050 62840 3056 62852
rect 3108 62840 3114 62892
rect 10134 62880 10140 62892
rect 10095 62852 10140 62880
rect 10134 62840 10140 62852
rect 10192 62840 10198 62892
rect 2314 62812 2320 62824
rect 2148 62784 2320 62812
rect 2314 62772 2320 62784
rect 2372 62772 2378 62824
rect 2685 62815 2743 62821
rect 2685 62781 2697 62815
rect 2731 62812 2743 62815
rect 3142 62812 3148 62824
rect 2731 62784 3148 62812
rect 2731 62781 2743 62784
rect 2685 62775 2743 62781
rect 3142 62772 3148 62784
rect 3200 62812 3206 62824
rect 3602 62812 3608 62824
rect 3200 62784 3608 62812
rect 3200 62772 3206 62784
rect 3602 62772 3608 62784
rect 3660 62772 3666 62824
rect 1673 62679 1731 62685
rect 1673 62645 1685 62679
rect 1719 62676 1731 62679
rect 8570 62676 8576 62688
rect 1719 62648 8576 62676
rect 1719 62645 1731 62648
rect 1673 62639 1731 62645
rect 8570 62636 8576 62648
rect 8628 62636 8634 62688
rect 1104 62586 10856 62608
rect 1104 62534 2582 62586
rect 2634 62534 2646 62586
rect 2698 62534 2710 62586
rect 2762 62534 2774 62586
rect 2826 62534 2838 62586
rect 2890 62534 5845 62586
rect 5897 62534 5909 62586
rect 5961 62534 5973 62586
rect 6025 62534 6037 62586
rect 6089 62534 6101 62586
rect 6153 62534 9109 62586
rect 9161 62534 9173 62586
rect 9225 62534 9237 62586
rect 9289 62534 9301 62586
rect 9353 62534 9365 62586
rect 9417 62534 10856 62586
rect 1104 62512 10856 62534
rect 2225 62407 2283 62413
rect 2225 62373 2237 62407
rect 2271 62404 2283 62407
rect 4614 62404 4620 62416
rect 2271 62376 4620 62404
rect 2271 62373 2283 62376
rect 2225 62367 2283 62373
rect 4614 62364 4620 62376
rect 4672 62364 4678 62416
rect 1673 62271 1731 62277
rect 1673 62237 1685 62271
rect 1719 62237 1731 62271
rect 1673 62231 1731 62237
rect 1394 62092 1400 62144
rect 1452 62132 1458 62144
rect 1489 62135 1547 62141
rect 1489 62132 1501 62135
rect 1452 62104 1501 62132
rect 1452 62092 1458 62104
rect 1489 62101 1501 62104
rect 1535 62101 1547 62135
rect 1688 62132 1716 62231
rect 2314 62228 2320 62280
rect 2372 62277 2378 62280
rect 2372 62271 2415 62277
rect 2403 62237 2415 62271
rect 2372 62231 2415 62237
rect 2777 62271 2835 62277
rect 2777 62237 2789 62271
rect 2823 62268 2835 62271
rect 3050 62268 3056 62280
rect 2823 62240 3056 62268
rect 2823 62237 2835 62240
rect 2777 62231 2835 62237
rect 2372 62228 2378 62231
rect 3050 62228 3056 62240
rect 3108 62228 3114 62280
rect 1946 62160 1952 62212
rect 2004 62200 2010 62212
rect 2501 62203 2559 62209
rect 2501 62200 2513 62203
rect 2004 62172 2513 62200
rect 2004 62160 2010 62172
rect 2501 62169 2513 62172
rect 2547 62169 2559 62203
rect 2501 62163 2559 62169
rect 2593 62203 2651 62209
rect 2593 62169 2605 62203
rect 2639 62200 2651 62203
rect 9950 62200 9956 62212
rect 2639 62172 9956 62200
rect 2639 62169 2651 62172
rect 2593 62163 2651 62169
rect 9950 62160 9956 62172
rect 10008 62160 10014 62212
rect 7282 62132 7288 62144
rect 1688 62104 7288 62132
rect 1489 62095 1547 62101
rect 7282 62092 7288 62104
rect 7340 62092 7346 62144
rect 1104 62042 10856 62064
rect 1104 61990 4213 62042
rect 4265 61990 4277 62042
rect 4329 61990 4341 62042
rect 4393 61990 4405 62042
rect 4457 61990 4469 62042
rect 4521 61990 7477 62042
rect 7529 61990 7541 62042
rect 7593 61990 7605 62042
rect 7657 61990 7669 62042
rect 7721 61990 7733 62042
rect 7785 61990 10856 62042
rect 1104 61968 10856 61990
rect 2222 61820 2228 61872
rect 2280 61860 2286 61872
rect 2501 61863 2559 61869
rect 2501 61860 2513 61863
rect 2280 61832 2513 61860
rect 2280 61820 2286 61832
rect 2501 61829 2513 61832
rect 2547 61829 2559 61863
rect 2501 61823 2559 61829
rect 290 61752 296 61804
rect 348 61792 354 61804
rect 1673 61795 1731 61801
rect 1673 61792 1685 61795
rect 348 61764 1685 61792
rect 348 61752 354 61764
rect 1673 61761 1685 61764
rect 1719 61761 1731 61795
rect 1673 61755 1731 61761
rect 2314 61752 2320 61804
rect 2372 61801 2378 61804
rect 2372 61795 2415 61801
rect 2403 61761 2415 61795
rect 2372 61755 2415 61761
rect 2593 61795 2651 61801
rect 2593 61761 2605 61795
rect 2639 61761 2651 61795
rect 2593 61755 2651 61761
rect 2777 61795 2835 61801
rect 2777 61761 2789 61795
rect 2823 61792 2835 61795
rect 3050 61792 3056 61804
rect 2823 61764 3056 61792
rect 2823 61761 2835 61764
rect 2777 61755 2835 61761
rect 2372 61752 2378 61755
rect 2608 61724 2636 61755
rect 3050 61752 3056 61764
rect 3108 61752 3114 61804
rect 10134 61792 10140 61804
rect 10095 61764 10140 61792
rect 10134 61752 10140 61764
rect 10192 61752 10198 61804
rect 2608 61696 2774 61724
rect 2746 61656 2774 61696
rect 9953 61659 10011 61665
rect 9953 61656 9965 61659
rect 2746 61628 9965 61656
rect 9953 61625 9965 61628
rect 9999 61625 10011 61659
rect 9953 61619 10011 61625
rect 1486 61588 1492 61600
rect 1447 61560 1492 61588
rect 1486 61548 1492 61560
rect 1544 61548 1550 61600
rect 2225 61591 2283 61597
rect 2225 61557 2237 61591
rect 2271 61588 2283 61591
rect 8662 61588 8668 61600
rect 2271 61560 8668 61588
rect 2271 61557 2283 61560
rect 2225 61551 2283 61557
rect 8662 61548 8668 61560
rect 8720 61548 8726 61600
rect 1104 61498 10856 61520
rect 1104 61446 2582 61498
rect 2634 61446 2646 61498
rect 2698 61446 2710 61498
rect 2762 61446 2774 61498
rect 2826 61446 2838 61498
rect 2890 61446 5845 61498
rect 5897 61446 5909 61498
rect 5961 61446 5973 61498
rect 6025 61446 6037 61498
rect 6089 61446 6101 61498
rect 6153 61446 9109 61498
rect 9161 61446 9173 61498
rect 9225 61446 9237 61498
rect 9289 61446 9301 61498
rect 9353 61446 9365 61498
rect 9417 61446 10856 61498
rect 1104 61424 10856 61446
rect 2222 61384 2228 61396
rect 2183 61356 2228 61384
rect 2222 61344 2228 61356
rect 2280 61344 2286 61396
rect 1673 61183 1731 61189
rect 1673 61149 1685 61183
rect 1719 61149 1731 61183
rect 1673 61143 1731 61149
rect 2409 61183 2467 61189
rect 2409 61149 2421 61183
rect 2455 61180 2467 61183
rect 4890 61180 4896 61192
rect 2455 61152 4896 61180
rect 2455 61149 2467 61152
rect 2409 61143 2467 61149
rect 1688 61112 1716 61143
rect 4890 61140 4896 61152
rect 4948 61140 4954 61192
rect 5626 61112 5632 61124
rect 1688 61084 5632 61112
rect 5626 61072 5632 61084
rect 5684 61072 5690 61124
rect 1394 61004 1400 61056
rect 1452 61044 1458 61056
rect 1489 61047 1547 61053
rect 1489 61044 1501 61047
rect 1452 61016 1501 61044
rect 1452 61004 1458 61016
rect 1489 61013 1501 61016
rect 1535 61013 1547 61047
rect 1489 61007 1547 61013
rect 1104 60954 10856 60976
rect 1104 60902 4213 60954
rect 4265 60902 4277 60954
rect 4329 60902 4341 60954
rect 4393 60902 4405 60954
rect 4457 60902 4469 60954
rect 4521 60902 7477 60954
rect 7529 60902 7541 60954
rect 7593 60902 7605 60954
rect 7657 60902 7669 60954
rect 7721 60902 7733 60954
rect 7785 60902 10856 60954
rect 1104 60880 10856 60902
rect 937 60843 995 60849
rect 937 60809 949 60843
rect 983 60840 995 60843
rect 1670 60840 1676 60852
rect 983 60812 1676 60840
rect 983 60809 995 60812
rect 937 60803 995 60809
rect 1670 60800 1676 60812
rect 1728 60800 1734 60852
rect 9950 60840 9956 60852
rect 9911 60812 9956 60840
rect 9950 60800 9956 60812
rect 10008 60800 10014 60852
rect 474 60664 480 60716
rect 532 60704 538 60716
rect 1673 60707 1731 60713
rect 1673 60704 1685 60707
rect 532 60676 1685 60704
rect 532 60664 538 60676
rect 1673 60673 1685 60676
rect 1719 60673 1731 60707
rect 10134 60704 10140 60716
rect 10095 60676 10140 60704
rect 1673 60667 1731 60673
rect 10134 60664 10140 60676
rect 10192 60664 10198 60716
rect 1486 60500 1492 60512
rect 1447 60472 1492 60500
rect 1486 60460 1492 60472
rect 1544 60460 1550 60512
rect 1104 60410 10856 60432
rect 1104 60358 2582 60410
rect 2634 60358 2646 60410
rect 2698 60358 2710 60410
rect 2762 60358 2774 60410
rect 2826 60358 2838 60410
rect 2890 60358 5845 60410
rect 5897 60358 5909 60410
rect 5961 60358 5973 60410
rect 6025 60358 6037 60410
rect 6089 60358 6101 60410
rect 6153 60358 9109 60410
rect 9161 60358 9173 60410
rect 9225 60358 9237 60410
rect 9289 60358 9301 60410
rect 9353 60358 9365 60410
rect 9417 60358 10856 60410
rect 1104 60336 10856 60358
rect 1673 60095 1731 60101
rect 1673 60061 1685 60095
rect 1719 60092 1731 60095
rect 6270 60092 6276 60104
rect 1719 60064 6276 60092
rect 1719 60061 1731 60064
rect 1673 60055 1731 60061
rect 6270 60052 6276 60064
rect 6328 60052 6334 60104
rect 1394 59916 1400 59968
rect 1452 59956 1458 59968
rect 1489 59959 1547 59965
rect 1489 59956 1501 59959
rect 1452 59928 1501 59956
rect 1452 59916 1458 59928
rect 1489 59925 1501 59928
rect 1535 59925 1547 59959
rect 1489 59919 1547 59925
rect 1104 59866 10856 59888
rect 1104 59814 4213 59866
rect 4265 59814 4277 59866
rect 4329 59814 4341 59866
rect 4393 59814 4405 59866
rect 4457 59814 4469 59866
rect 4521 59814 7477 59866
rect 7529 59814 7541 59866
rect 7593 59814 7605 59866
rect 7657 59814 7669 59866
rect 7721 59814 7733 59866
rect 7785 59814 10856 59866
rect 1104 59792 10856 59814
rect 566 59576 572 59628
rect 624 59616 630 59628
rect 1673 59619 1731 59625
rect 1673 59616 1685 59619
rect 624 59588 1685 59616
rect 624 59576 630 59588
rect 1673 59585 1685 59588
rect 1719 59585 1731 59619
rect 1673 59579 1731 59585
rect 2409 59619 2467 59625
rect 2409 59585 2421 59619
rect 2455 59616 2467 59619
rect 5350 59616 5356 59628
rect 2455 59588 5356 59616
rect 2455 59585 2467 59588
rect 2409 59579 2467 59585
rect 5350 59576 5356 59588
rect 5408 59576 5414 59628
rect 10134 59616 10140 59628
rect 10095 59588 10140 59616
rect 10134 59576 10140 59588
rect 10192 59576 10198 59628
rect 2222 59480 2228 59492
rect 2183 59452 2228 59480
rect 2222 59440 2228 59452
rect 2280 59440 2286 59492
rect 1486 59412 1492 59424
rect 1447 59384 1492 59412
rect 1486 59372 1492 59384
rect 1544 59372 1550 59424
rect 9950 59412 9956 59424
rect 9911 59384 9956 59412
rect 9950 59372 9956 59384
rect 10008 59372 10014 59424
rect 1104 59322 10856 59344
rect 1104 59270 2582 59322
rect 2634 59270 2646 59322
rect 2698 59270 2710 59322
rect 2762 59270 2774 59322
rect 2826 59270 2838 59322
rect 2890 59270 5845 59322
rect 5897 59270 5909 59322
rect 5961 59270 5973 59322
rect 6025 59270 6037 59322
rect 6089 59270 6101 59322
rect 6153 59270 9109 59322
rect 9161 59270 9173 59322
rect 9225 59270 9237 59322
rect 9289 59270 9301 59322
rect 9353 59270 9365 59322
rect 9417 59270 10856 59322
rect 1104 59248 10856 59270
rect 1397 59143 1455 59149
rect 1397 59109 1409 59143
rect 1443 59140 1455 59143
rect 3878 59140 3884 59152
rect 1443 59112 3884 59140
rect 1443 59109 1455 59112
rect 1397 59103 1455 59109
rect 3878 59100 3884 59112
rect 3936 59100 3942 59152
rect 2314 59072 2320 59084
rect 1688 59044 2320 59072
rect 1688 59013 1716 59044
rect 2314 59032 2320 59044
rect 2372 59032 2378 59084
rect 1581 59007 1639 59013
rect 1581 59004 1593 59007
rect 1412 58976 1593 59004
rect 1412 58880 1440 58976
rect 1581 58973 1593 58976
rect 1627 58973 1639 59007
rect 1581 58967 1639 58973
rect 1673 59007 1731 59013
rect 1673 58973 1685 59007
rect 1719 58973 1731 59007
rect 1673 58967 1731 58973
rect 1949 59007 2007 59013
rect 1949 58973 1961 59007
rect 1995 59004 2007 59007
rect 2222 59004 2228 59016
rect 1995 58976 2228 59004
rect 1995 58973 2007 58976
rect 1949 58967 2007 58973
rect 2222 58964 2228 58976
rect 2280 58964 2286 59016
rect 2685 59007 2743 59013
rect 2685 58973 2697 59007
rect 2731 59004 2743 59007
rect 5442 59004 5448 59016
rect 2731 58976 5448 59004
rect 2731 58973 2743 58976
rect 2685 58967 2743 58973
rect 5442 58964 5448 58976
rect 5500 58964 5506 59016
rect 1765 58939 1823 58945
rect 1765 58905 1777 58939
rect 1811 58936 1823 58939
rect 9950 58936 9956 58948
rect 1811 58908 9956 58936
rect 1811 58905 1823 58908
rect 1765 58899 1823 58905
rect 9950 58896 9956 58908
rect 10008 58896 10014 58948
rect 1394 58828 1400 58880
rect 1452 58828 1458 58880
rect 2501 58871 2559 58877
rect 2501 58837 2513 58871
rect 2547 58868 2559 58871
rect 2774 58868 2780 58880
rect 2547 58840 2780 58868
rect 2547 58837 2559 58840
rect 2501 58831 2559 58837
rect 2774 58828 2780 58840
rect 2832 58828 2838 58880
rect 1104 58778 10856 58800
rect 1104 58726 4213 58778
rect 4265 58726 4277 58778
rect 4329 58726 4341 58778
rect 4393 58726 4405 58778
rect 4457 58726 4469 58778
rect 4521 58726 7477 58778
rect 7529 58726 7541 58778
rect 7593 58726 7605 58778
rect 7657 58726 7669 58778
rect 7721 58726 7733 58778
rect 7785 58726 10856 58778
rect 1104 58704 10856 58726
rect 1762 58624 1768 58676
rect 1820 58624 1826 58676
rect 1673 58599 1731 58605
rect 1673 58565 1685 58599
rect 1719 58596 1731 58599
rect 1780 58596 1808 58624
rect 1719 58568 1808 58596
rect 1719 58565 1731 58568
rect 1673 58559 1731 58565
rect 1394 58488 1400 58540
rect 1452 58528 1458 58540
rect 1581 58531 1639 58537
rect 1581 58528 1593 58531
rect 1452 58500 1593 58528
rect 1452 58488 1458 58500
rect 1581 58497 1593 58500
rect 1627 58497 1639 58531
rect 1581 58491 1639 58497
rect 1765 58531 1823 58537
rect 1765 58497 1777 58531
rect 1811 58497 1823 58531
rect 1765 58491 1823 58497
rect 1949 58531 2007 58537
rect 1949 58497 1961 58531
rect 1995 58528 2007 58531
rect 2222 58528 2228 58540
rect 1995 58500 2228 58528
rect 1995 58497 2007 58500
rect 1949 58491 2007 58497
rect 1780 58460 1808 58491
rect 2222 58488 2228 58500
rect 2280 58488 2286 58540
rect 2685 58531 2743 58537
rect 2685 58497 2697 58531
rect 2731 58528 2743 58531
rect 4798 58528 4804 58540
rect 2731 58500 4804 58528
rect 2731 58497 2743 58500
rect 2685 58491 2743 58497
rect 4798 58488 4804 58500
rect 4856 58488 4862 58540
rect 10134 58528 10140 58540
rect 10095 58500 10140 58528
rect 10134 58488 10140 58500
rect 10192 58488 10198 58540
rect 1780 58432 2774 58460
rect 2746 58392 2774 58432
rect 9953 58395 10011 58401
rect 9953 58392 9965 58395
rect 2746 58364 9965 58392
rect 9953 58361 9965 58364
rect 9999 58361 10011 58395
rect 9953 58355 10011 58361
rect 1397 58327 1455 58333
rect 1397 58293 1409 58327
rect 1443 58324 1455 58327
rect 1578 58324 1584 58336
rect 1443 58296 1584 58324
rect 1443 58293 1455 58296
rect 1397 58287 1455 58293
rect 1578 58284 1584 58296
rect 1636 58284 1642 58336
rect 2498 58324 2504 58336
rect 2459 58296 2504 58324
rect 2498 58284 2504 58296
rect 2556 58284 2562 58336
rect 1104 58234 10856 58256
rect 1104 58182 2582 58234
rect 2634 58182 2646 58234
rect 2698 58182 2710 58234
rect 2762 58182 2774 58234
rect 2826 58182 2838 58234
rect 2890 58182 5845 58234
rect 5897 58182 5909 58234
rect 5961 58182 5973 58234
rect 6025 58182 6037 58234
rect 6089 58182 6101 58234
rect 6153 58182 9109 58234
rect 9161 58182 9173 58234
rect 9225 58182 9237 58234
rect 9289 58182 9301 58234
rect 9353 58182 9365 58234
rect 9417 58182 10856 58234
rect 1104 58160 10856 58182
rect 2130 58012 2136 58064
rect 2188 58052 2194 58064
rect 2590 58052 2596 58064
rect 2188 58024 2596 58052
rect 2188 58012 2194 58024
rect 2590 58012 2596 58024
rect 2648 58012 2654 58064
rect 1486 57944 1492 57996
rect 1544 57984 1550 57996
rect 1544 57956 1808 57984
rect 1544 57944 1550 57956
rect 1394 57916 1400 57928
rect 1355 57888 1400 57916
rect 1394 57876 1400 57888
rect 1452 57876 1458 57928
rect 1670 57916 1676 57928
rect 1631 57888 1676 57916
rect 1670 57876 1676 57888
rect 1728 57876 1734 57928
rect 1780 57925 1808 57956
rect 2038 57944 2044 57996
rect 2096 57984 2102 57996
rect 2314 57984 2320 57996
rect 2096 57956 2320 57984
rect 2096 57944 2102 57956
rect 2314 57944 2320 57956
rect 2372 57944 2378 57996
rect 2608 57956 2820 57984
rect 1765 57919 1823 57925
rect 1765 57885 1777 57919
rect 1811 57916 1823 57919
rect 2409 57919 2467 57925
rect 1811 57888 2268 57916
rect 1811 57885 1823 57888
rect 1765 57879 1823 57885
rect 1581 57851 1639 57857
rect 1581 57817 1593 57851
rect 1627 57848 1639 57851
rect 2130 57848 2136 57860
rect 1627 57820 2136 57848
rect 1627 57817 1639 57820
rect 1581 57811 1639 57817
rect 2130 57808 2136 57820
rect 2188 57808 2194 57860
rect 2240 57848 2268 57888
rect 2409 57885 2421 57919
rect 2455 57916 2467 57919
rect 2608 57916 2636 57956
rect 2455 57888 2636 57916
rect 2685 57919 2743 57925
rect 2455 57885 2467 57888
rect 2409 57879 2467 57885
rect 2685 57885 2697 57919
rect 2731 57885 2743 57919
rect 2792 57916 2820 57956
rect 3510 57916 3516 57928
rect 2792 57888 3516 57916
rect 2685 57879 2743 57885
rect 2700 57848 2728 57879
rect 3510 57876 3516 57888
rect 3568 57876 3574 57928
rect 2240 57820 2728 57848
rect 1949 57783 2007 57789
rect 1949 57749 1961 57783
rect 1995 57780 2007 57783
rect 2038 57780 2044 57792
rect 1995 57752 2044 57780
rect 1995 57749 2007 57752
rect 1949 57743 2007 57749
rect 2038 57740 2044 57752
rect 2096 57740 2102 57792
rect 1104 57690 10856 57712
rect 1104 57638 4213 57690
rect 4265 57638 4277 57690
rect 4329 57638 4341 57690
rect 4393 57638 4405 57690
rect 4457 57638 4469 57690
rect 4521 57638 7477 57690
rect 7529 57638 7541 57690
rect 7593 57638 7605 57690
rect 7657 57638 7669 57690
rect 7721 57638 7733 57690
rect 7785 57638 10856 57690
rect 1104 57616 10856 57638
rect 1394 57576 1400 57588
rect 1307 57548 1400 57576
rect 1394 57536 1400 57548
rect 1452 57576 1458 57588
rect 2222 57576 2228 57588
rect 1452 57548 2228 57576
rect 1452 57536 1458 57548
rect 2222 57536 2228 57548
rect 2280 57536 2286 57588
rect 1412 57449 1440 57536
rect 1581 57511 1639 57517
rect 1581 57477 1593 57511
rect 1627 57508 1639 57511
rect 9858 57508 9864 57520
rect 1627 57480 9864 57508
rect 1627 57477 1639 57480
rect 1581 57471 1639 57477
rect 9858 57468 9864 57480
rect 9916 57468 9922 57520
rect 1397 57443 1455 57449
rect 1397 57409 1409 57443
rect 1443 57409 1455 57443
rect 1670 57440 1676 57452
rect 1631 57412 1676 57440
rect 1397 57403 1455 57409
rect 1670 57400 1676 57412
rect 1728 57400 1734 57452
rect 1765 57443 1823 57449
rect 1765 57409 1777 57443
rect 1811 57409 1823 57443
rect 1765 57403 1823 57409
rect 1486 57332 1492 57384
rect 1544 57372 1550 57384
rect 1780 57372 1808 57403
rect 2222 57400 2228 57452
rect 2280 57440 2286 57452
rect 2685 57443 2743 57449
rect 2685 57440 2697 57443
rect 2280 57412 2697 57440
rect 2280 57400 2286 57412
rect 2685 57409 2697 57412
rect 2731 57409 2743 57443
rect 2685 57403 2743 57409
rect 3697 57443 3755 57449
rect 3697 57409 3709 57443
rect 3743 57440 3755 57443
rect 6178 57440 6184 57452
rect 3743 57412 6184 57440
rect 3743 57409 3755 57412
rect 3697 57403 3755 57409
rect 6178 57400 6184 57412
rect 6236 57400 6242 57452
rect 10134 57440 10140 57452
rect 10095 57412 10140 57440
rect 10134 57400 10140 57412
rect 10192 57400 10198 57452
rect 1544 57344 1808 57372
rect 2409 57375 2467 57381
rect 1544 57332 1550 57344
rect 2409 57341 2421 57375
rect 2455 57372 2467 57375
rect 3050 57372 3056 57384
rect 2455 57344 3056 57372
rect 2455 57341 2467 57344
rect 2409 57335 2467 57341
rect 1394 57264 1400 57316
rect 1452 57304 1458 57316
rect 2424 57304 2452 57335
rect 3050 57332 3056 57344
rect 3108 57332 3114 57384
rect 1452 57276 2452 57304
rect 1452 57264 1458 57276
rect 3142 57264 3148 57316
rect 3200 57304 3206 57316
rect 3881 57307 3939 57313
rect 3881 57304 3893 57307
rect 3200 57276 3893 57304
rect 3200 57264 3206 57276
rect 3881 57273 3893 57276
rect 3927 57273 3939 57307
rect 3881 57267 3939 57273
rect 1949 57239 2007 57245
rect 1949 57205 1961 57239
rect 1995 57236 2007 57239
rect 3694 57236 3700 57248
rect 1995 57208 3700 57236
rect 1995 57205 2007 57208
rect 1949 57199 2007 57205
rect 3694 57196 3700 57208
rect 3752 57196 3758 57248
rect 9950 57236 9956 57248
rect 9911 57208 9956 57236
rect 9950 57196 9956 57208
rect 10008 57196 10014 57248
rect 1104 57146 10856 57168
rect 1104 57094 2582 57146
rect 2634 57094 2646 57146
rect 2698 57094 2710 57146
rect 2762 57094 2774 57146
rect 2826 57094 2838 57146
rect 2890 57094 5845 57146
rect 5897 57094 5909 57146
rect 5961 57094 5973 57146
rect 6025 57094 6037 57146
rect 6089 57094 6101 57146
rect 6153 57094 9109 57146
rect 9161 57094 9173 57146
rect 9225 57094 9237 57146
rect 9289 57094 9301 57146
rect 9353 57094 9365 57146
rect 9417 57094 10856 57146
rect 1104 57072 10856 57094
rect 1670 56992 1676 57044
rect 1728 57032 1734 57044
rect 1946 57032 1952 57044
rect 1728 57004 1952 57032
rect 1728 56992 1734 57004
rect 1946 56992 1952 57004
rect 2004 56992 2010 57044
rect 2130 56992 2136 57044
rect 2188 57032 2194 57044
rect 9950 57032 9956 57044
rect 2188 57004 9956 57032
rect 2188 56992 2194 57004
rect 9950 56992 9956 57004
rect 10008 56992 10014 57044
rect 750 56856 756 56908
rect 808 56896 814 56908
rect 1670 56896 1676 56908
rect 808 56868 1676 56896
rect 808 56856 814 56868
rect 1670 56856 1676 56868
rect 1728 56856 1734 56908
rect 1486 56788 1492 56840
rect 1544 56828 1550 56840
rect 1581 56831 1639 56837
rect 1581 56828 1593 56831
rect 1544 56800 1593 56828
rect 1544 56788 1550 56800
rect 1581 56797 1593 56800
rect 1627 56797 1639 56831
rect 1854 56828 1860 56840
rect 1581 56791 1639 56797
rect 1688 56800 1860 56828
rect 1688 56769 1716 56800
rect 1854 56788 1860 56800
rect 1912 56788 1918 56840
rect 1949 56831 2007 56837
rect 1949 56797 1961 56831
rect 1995 56828 2007 56831
rect 2222 56828 2228 56840
rect 1995 56800 2228 56828
rect 1995 56797 2007 56800
rect 1949 56791 2007 56797
rect 2222 56788 2228 56800
rect 2280 56788 2286 56840
rect 2685 56831 2743 56837
rect 2685 56797 2697 56831
rect 2731 56828 2743 56831
rect 6362 56828 6368 56840
rect 2731 56800 6368 56828
rect 2731 56797 2743 56800
rect 2685 56791 2743 56797
rect 6362 56788 6368 56800
rect 6420 56788 6426 56840
rect 1673 56763 1731 56769
rect 1673 56729 1685 56763
rect 1719 56729 1731 56763
rect 1673 56723 1731 56729
rect 1765 56763 1823 56769
rect 1765 56729 1777 56763
rect 1811 56760 1823 56763
rect 9950 56760 9956 56772
rect 1811 56732 9956 56760
rect 1811 56729 1823 56732
rect 1765 56723 1823 56729
rect 9950 56720 9956 56732
rect 10008 56720 10014 56772
rect 658 56652 664 56704
rect 716 56692 722 56704
rect 1302 56692 1308 56704
rect 716 56664 1308 56692
rect 716 56652 722 56664
rect 1302 56652 1308 56664
rect 1360 56652 1366 56704
rect 1397 56695 1455 56701
rect 1397 56661 1409 56695
rect 1443 56692 1455 56695
rect 1946 56692 1952 56704
rect 1443 56664 1952 56692
rect 1443 56661 1455 56664
rect 1397 56655 1455 56661
rect 1946 56652 1952 56664
rect 2004 56652 2010 56704
rect 2498 56692 2504 56704
rect 2459 56664 2504 56692
rect 2498 56652 2504 56664
rect 2556 56652 2562 56704
rect 3050 56652 3056 56704
rect 3108 56692 3114 56704
rect 4706 56692 4712 56704
rect 3108 56664 4712 56692
rect 3108 56652 3114 56664
rect 4706 56652 4712 56664
rect 4764 56652 4770 56704
rect 1104 56602 10856 56624
rect 1104 56550 4213 56602
rect 4265 56550 4277 56602
rect 4329 56550 4341 56602
rect 4393 56550 4405 56602
rect 4457 56550 4469 56602
rect 4521 56550 7477 56602
rect 7529 56550 7541 56602
rect 7593 56550 7605 56602
rect 7657 56550 7669 56602
rect 7721 56550 7733 56602
rect 7785 56550 10856 56602
rect 1104 56528 10856 56550
rect 1394 56448 1400 56500
rect 1452 56488 1458 56500
rect 1854 56488 1860 56500
rect 1452 56460 1860 56488
rect 1452 56448 1458 56460
rect 1854 56448 1860 56460
rect 1912 56448 1918 56500
rect 3053 56491 3111 56497
rect 3053 56457 3065 56491
rect 3099 56488 3111 56491
rect 3510 56488 3516 56500
rect 3099 56460 3516 56488
rect 3099 56457 3111 56460
rect 3053 56451 3111 56457
rect 3510 56448 3516 56460
rect 3568 56448 3574 56500
rect 9950 56488 9956 56500
rect 9911 56460 9956 56488
rect 9950 56448 9956 56460
rect 10008 56448 10014 56500
rect 1394 56312 1400 56364
rect 1452 56352 1458 56364
rect 1673 56355 1731 56361
rect 1673 56352 1685 56355
rect 1452 56324 1685 56352
rect 1452 56312 1458 56324
rect 1673 56321 1685 56324
rect 1719 56321 1731 56355
rect 1673 56315 1731 56321
rect 2133 56355 2191 56361
rect 2133 56321 2145 56355
rect 2179 56352 2191 56355
rect 2961 56355 3019 56361
rect 2179 56324 2774 56352
rect 2179 56321 2191 56324
rect 2133 56315 2191 56321
rect 2746 56284 2774 56324
rect 2961 56321 2973 56355
rect 3007 56352 3019 56355
rect 3142 56352 3148 56364
rect 3007 56324 3148 56352
rect 3007 56321 3019 56324
rect 2961 56315 3019 56321
rect 3142 56312 3148 56324
rect 3200 56312 3206 56364
rect 10134 56352 10140 56364
rect 10095 56324 10140 56352
rect 10134 56312 10140 56324
rect 10192 56312 10198 56364
rect 6546 56284 6552 56296
rect 2746 56256 6552 56284
rect 6546 56244 6552 56256
rect 6604 56244 6610 56296
rect 2314 56216 2320 56228
rect 2275 56188 2320 56216
rect 2314 56176 2320 56188
rect 2372 56176 2378 56228
rect 1486 56148 1492 56160
rect 1447 56120 1492 56148
rect 1486 56108 1492 56120
rect 1544 56108 1550 56160
rect 1104 56058 10856 56080
rect 1104 56006 2582 56058
rect 2634 56006 2646 56058
rect 2698 56006 2710 56058
rect 2762 56006 2774 56058
rect 2826 56006 2838 56058
rect 2890 56006 5845 56058
rect 5897 56006 5909 56058
rect 5961 56006 5973 56058
rect 6025 56006 6037 56058
rect 6089 56006 6101 56058
rect 6153 56006 9109 56058
rect 9161 56006 9173 56058
rect 9225 56006 9237 56058
rect 9289 56006 9301 56058
rect 9353 56006 9365 56058
rect 9417 56006 10856 56058
rect 1104 55984 10856 56006
rect 3050 55904 3056 55956
rect 3108 55944 3114 55956
rect 3418 55944 3424 55956
rect 3108 55916 3424 55944
rect 3108 55904 3114 55916
rect 3418 55904 3424 55916
rect 3476 55904 3482 55956
rect 1673 55743 1731 55749
rect 1673 55709 1685 55743
rect 1719 55740 1731 55743
rect 1719 55712 4752 55740
rect 1719 55709 1731 55712
rect 1673 55703 1731 55709
rect 4724 55616 4752 55712
rect 1486 55604 1492 55616
rect 1447 55576 1492 55604
rect 1486 55564 1492 55576
rect 1544 55564 1550 55616
rect 3142 55564 3148 55616
rect 3200 55604 3206 55616
rect 3694 55604 3700 55616
rect 3200 55576 3700 55604
rect 3200 55564 3206 55576
rect 3694 55564 3700 55576
rect 3752 55564 3758 55616
rect 4706 55564 4712 55616
rect 4764 55564 4770 55616
rect 1104 55514 10856 55536
rect 1104 55462 4213 55514
rect 4265 55462 4277 55514
rect 4329 55462 4341 55514
rect 4393 55462 4405 55514
rect 4457 55462 4469 55514
rect 4521 55462 7477 55514
rect 7529 55462 7541 55514
rect 7593 55462 7605 55514
rect 7657 55462 7669 55514
rect 7721 55462 7733 55514
rect 7785 55462 10856 55514
rect 1104 55440 10856 55462
rect 2958 55360 2964 55412
rect 3016 55400 3022 55412
rect 3602 55400 3608 55412
rect 3016 55372 3608 55400
rect 3016 55360 3022 55372
rect 3602 55360 3608 55372
rect 3660 55360 3666 55412
rect 9858 55360 9864 55412
rect 9916 55400 9922 55412
rect 9953 55403 10011 55409
rect 9953 55400 9965 55403
rect 9916 55372 9965 55400
rect 9916 55360 9922 55372
rect 9953 55369 9965 55372
rect 9999 55369 10011 55403
rect 9953 55363 10011 55369
rect 7834 55332 7840 55344
rect 1688 55304 7840 55332
rect 1688 55273 1716 55304
rect 7834 55292 7840 55304
rect 7892 55292 7898 55344
rect 1673 55267 1731 55273
rect 1673 55233 1685 55267
rect 1719 55233 1731 55267
rect 1673 55227 1731 55233
rect 2409 55267 2467 55273
rect 2409 55233 2421 55267
rect 2455 55264 2467 55267
rect 3142 55264 3148 55276
rect 2455 55236 3148 55264
rect 2455 55233 2467 55236
rect 2409 55227 2467 55233
rect 3142 55224 3148 55236
rect 3200 55224 3206 55276
rect 10134 55264 10140 55276
rect 10095 55236 10140 55264
rect 10134 55224 10140 55236
rect 10192 55224 10198 55276
rect 1486 55060 1492 55072
rect 1447 55032 1492 55060
rect 1486 55020 1492 55032
rect 1544 55020 1550 55072
rect 2222 55060 2228 55072
rect 2183 55032 2228 55060
rect 2222 55020 2228 55032
rect 2280 55020 2286 55072
rect 1104 54970 10856 54992
rect 1104 54918 2582 54970
rect 2634 54918 2646 54970
rect 2698 54918 2710 54970
rect 2762 54918 2774 54970
rect 2826 54918 2838 54970
rect 2890 54918 5845 54970
rect 5897 54918 5909 54970
rect 5961 54918 5973 54970
rect 6025 54918 6037 54970
rect 6089 54918 6101 54970
rect 6153 54918 9109 54970
rect 9161 54918 9173 54970
rect 9225 54918 9237 54970
rect 9289 54918 9301 54970
rect 9353 54918 9365 54970
rect 9417 54918 10856 54970
rect 1104 54896 10856 54918
rect 3878 54816 3884 54868
rect 3936 54856 3942 54868
rect 3936 54828 4016 54856
rect 3936 54816 3942 54828
rect 3988 54664 4016 54828
rect 658 54612 664 54664
rect 716 54652 722 54664
rect 1673 54655 1731 54661
rect 1673 54652 1685 54655
rect 716 54624 1685 54652
rect 716 54612 722 54624
rect 1673 54621 1685 54624
rect 1719 54621 1731 54655
rect 1673 54615 1731 54621
rect 3970 54612 3976 54664
rect 4028 54612 4034 54664
rect 1394 54476 1400 54528
rect 1452 54516 1458 54528
rect 1489 54519 1547 54525
rect 1489 54516 1501 54519
rect 1452 54488 1501 54516
rect 1452 54476 1458 54488
rect 1489 54485 1501 54488
rect 1535 54485 1547 54519
rect 1489 54479 1547 54485
rect 1104 54426 10856 54448
rect 1104 54374 4213 54426
rect 4265 54374 4277 54426
rect 4329 54374 4341 54426
rect 4393 54374 4405 54426
rect 4457 54374 4469 54426
rect 4521 54374 7477 54426
rect 7529 54374 7541 54426
rect 7593 54374 7605 54426
rect 7657 54374 7669 54426
rect 7721 54374 7733 54426
rect 7785 54374 10856 54426
rect 1104 54352 10856 54374
rect 1673 54179 1731 54185
rect 1673 54145 1685 54179
rect 1719 54145 1731 54179
rect 1673 54139 1731 54145
rect 2409 54179 2467 54185
rect 2409 54145 2421 54179
rect 2455 54176 2467 54179
rect 7006 54176 7012 54188
rect 2455 54148 7012 54176
rect 2455 54145 2467 54148
rect 2409 54139 2467 54145
rect 1688 54108 1716 54139
rect 7006 54136 7012 54148
rect 7064 54136 7070 54188
rect 10134 54176 10140 54188
rect 10095 54148 10140 54176
rect 10134 54136 10140 54148
rect 10192 54136 10198 54188
rect 7098 54108 7104 54120
rect 1688 54080 7104 54108
rect 7098 54068 7104 54080
rect 7156 54068 7162 54120
rect 2222 54040 2228 54052
rect 2183 54012 2228 54040
rect 2222 54000 2228 54012
rect 2280 54000 2286 54052
rect 1486 53972 1492 53984
rect 1447 53944 1492 53972
rect 1486 53932 1492 53944
rect 1544 53932 1550 53984
rect 9950 53972 9956 53984
rect 9911 53944 9956 53972
rect 9950 53932 9956 53944
rect 10008 53932 10014 53984
rect 1104 53882 10856 53904
rect 1104 53830 2582 53882
rect 2634 53830 2646 53882
rect 2698 53830 2710 53882
rect 2762 53830 2774 53882
rect 2826 53830 2838 53882
rect 2890 53830 5845 53882
rect 5897 53830 5909 53882
rect 5961 53830 5973 53882
rect 6025 53830 6037 53882
rect 6089 53830 6101 53882
rect 6153 53830 9109 53882
rect 9161 53830 9173 53882
rect 9225 53830 9237 53882
rect 9289 53830 9301 53882
rect 9353 53830 9365 53882
rect 9417 53830 10856 53882
rect 1104 53808 10856 53830
rect 1210 53728 1216 53780
rect 1268 53768 1274 53780
rect 1854 53768 1860 53780
rect 1268 53740 1860 53768
rect 1268 53728 1274 53740
rect 1854 53728 1860 53740
rect 1912 53728 1918 53780
rect 2038 53728 2044 53780
rect 2096 53768 2102 53780
rect 2498 53768 2504 53780
rect 2096 53740 2504 53768
rect 2096 53728 2102 53740
rect 2498 53728 2504 53740
rect 2556 53728 2562 53780
rect 2869 53771 2927 53777
rect 2869 53737 2881 53771
rect 2915 53768 2927 53771
rect 4062 53768 4068 53780
rect 2915 53740 4068 53768
rect 2915 53737 2927 53740
rect 2869 53731 2927 53737
rect 4062 53728 4068 53740
rect 4120 53728 4126 53780
rect 2498 53592 2504 53644
rect 2556 53632 2562 53644
rect 2958 53632 2964 53644
rect 2556 53604 2964 53632
rect 2556 53592 2562 53604
rect 2958 53592 2964 53604
rect 3016 53592 3022 53644
rect 753 53567 811 53573
rect 753 53533 765 53567
rect 799 53564 811 53567
rect 1673 53567 1731 53573
rect 1673 53564 1685 53567
rect 799 53536 1685 53564
rect 799 53533 811 53536
rect 753 53527 811 53533
rect 1673 53533 1685 53536
rect 1719 53533 1731 53567
rect 1673 53527 1731 53533
rect 2133 53567 2191 53573
rect 2133 53533 2145 53567
rect 2179 53564 2191 53567
rect 2179 53536 2774 53564
rect 2179 53533 2191 53536
rect 2133 53527 2191 53533
rect 2746 53496 2774 53536
rect 2866 53524 2872 53576
rect 2924 53564 2930 53576
rect 3053 53567 3111 53573
rect 2924 53536 2969 53564
rect 2924 53524 2930 53536
rect 3053 53533 3065 53567
rect 3099 53564 3111 53567
rect 5442 53564 5448 53576
rect 3099 53536 5448 53564
rect 3099 53533 3111 53536
rect 3053 53527 3111 53533
rect 5442 53524 5448 53536
rect 5500 53524 5506 53576
rect 7190 53496 7196 53508
rect 2746 53468 7196 53496
rect 7190 53456 7196 53468
rect 7248 53456 7254 53508
rect 1394 53388 1400 53440
rect 1452 53428 1458 53440
rect 1489 53431 1547 53437
rect 1489 53428 1501 53431
rect 1452 53400 1501 53428
rect 1452 53388 1458 53400
rect 1489 53397 1501 53400
rect 1535 53397 1547 53431
rect 2314 53428 2320 53440
rect 2275 53400 2320 53428
rect 1489 53391 1547 53397
rect 2314 53388 2320 53400
rect 2372 53388 2378 53440
rect 1104 53338 10856 53360
rect 1104 53286 4213 53338
rect 4265 53286 4277 53338
rect 4329 53286 4341 53338
rect 4393 53286 4405 53338
rect 4457 53286 4469 53338
rect 4521 53286 7477 53338
rect 7529 53286 7541 53338
rect 7593 53286 7605 53338
rect 7657 53286 7669 53338
rect 7721 53286 7733 53338
rect 7785 53286 10856 53338
rect 1104 53264 10856 53286
rect 1946 53224 1952 53236
rect 1412 53196 1952 53224
rect 1412 53097 1440 53196
rect 1946 53184 1952 53196
rect 2004 53184 2010 53236
rect 3237 53227 3295 53233
rect 3237 53193 3249 53227
rect 3283 53224 3295 53227
rect 3326 53224 3332 53236
rect 3283 53196 3332 53224
rect 3283 53193 3295 53196
rect 3237 53187 3295 53193
rect 3326 53184 3332 53196
rect 3384 53184 3390 53236
rect 4062 53184 4068 53236
rect 4120 53224 4126 53236
rect 5258 53224 5264 53236
rect 4120 53196 5264 53224
rect 4120 53184 4126 53196
rect 5258 53184 5264 53196
rect 5316 53184 5322 53236
rect 1581 53159 1639 53165
rect 1581 53125 1593 53159
rect 1627 53156 1639 53159
rect 9950 53156 9956 53168
rect 1627 53128 9956 53156
rect 1627 53125 1639 53128
rect 1581 53119 1639 53125
rect 9950 53116 9956 53128
rect 10008 53116 10014 53168
rect 1397 53091 1455 53097
rect 1397 53057 1409 53091
rect 1443 53057 1455 53091
rect 1397 53051 1455 53057
rect 1673 53091 1731 53097
rect 1673 53057 1685 53091
rect 1719 53057 1731 53091
rect 1673 53051 1731 53057
rect 1765 53091 1823 53097
rect 1765 53057 1777 53091
rect 1811 53088 1823 53091
rect 1854 53088 1860 53100
rect 1811 53060 1860 53088
rect 1811 53057 1823 53060
rect 1765 53051 1823 53057
rect 1688 53020 1716 53051
rect 1854 53048 1860 53060
rect 1912 53048 1918 53100
rect 2685 53091 2743 53097
rect 2685 53057 2697 53091
rect 2731 53088 2743 53091
rect 3050 53088 3056 53100
rect 2731 53060 3056 53088
rect 2731 53057 2743 53060
rect 2685 53051 2743 53057
rect 3050 53048 3056 53060
rect 3108 53048 3114 53100
rect 3145 53091 3203 53097
rect 3145 53057 3157 53091
rect 3191 53057 3203 53091
rect 3326 53088 3332 53100
rect 3287 53060 3332 53088
rect 3145 53051 3203 53057
rect 2038 53020 2044 53032
rect 1688 52992 2044 53020
rect 2038 52980 2044 52992
rect 2096 52980 2102 53032
rect 3160 53020 3188 53051
rect 3326 53048 3332 53060
rect 3384 53048 3390 53100
rect 4614 53048 4620 53100
rect 4672 53088 4678 53100
rect 5258 53088 5264 53100
rect 4672 53060 5264 53088
rect 4672 53048 4678 53060
rect 5258 53048 5264 53060
rect 5316 53048 5322 53100
rect 10134 53088 10140 53100
rect 10095 53060 10140 53088
rect 10134 53048 10140 53060
rect 10192 53048 10198 53100
rect 3160 52992 5396 53020
rect 5368 52964 5396 52992
rect 2866 52912 2872 52964
rect 2924 52952 2930 52964
rect 2924 52924 3096 52952
rect 2924 52912 2930 52924
rect 1949 52887 2007 52893
rect 1949 52853 1961 52887
rect 1995 52884 2007 52887
rect 2038 52884 2044 52896
rect 1995 52856 2044 52884
rect 1995 52853 2007 52856
rect 1949 52847 2007 52853
rect 2038 52844 2044 52856
rect 2096 52844 2102 52896
rect 2501 52887 2559 52893
rect 2501 52853 2513 52887
rect 2547 52884 2559 52887
rect 2958 52884 2964 52896
rect 2547 52856 2964 52884
rect 2547 52853 2559 52856
rect 2501 52847 2559 52853
rect 2958 52844 2964 52856
rect 3016 52844 3022 52896
rect 3068 52884 3096 52924
rect 5350 52912 5356 52964
rect 5408 52912 5414 52964
rect 3326 52884 3332 52896
rect 3068 52856 3332 52884
rect 3326 52844 3332 52856
rect 3384 52844 3390 52896
rect 9950 52884 9956 52896
rect 9911 52856 9956 52884
rect 9950 52844 9956 52856
rect 10008 52844 10014 52896
rect 1104 52794 10856 52816
rect 1104 52742 2582 52794
rect 2634 52742 2646 52794
rect 2698 52742 2710 52794
rect 2762 52742 2774 52794
rect 2826 52742 2838 52794
rect 2890 52742 5845 52794
rect 5897 52742 5909 52794
rect 5961 52742 5973 52794
rect 6025 52742 6037 52794
rect 6089 52742 6101 52794
rect 6153 52742 9109 52794
rect 9161 52742 9173 52794
rect 9225 52742 9237 52794
rect 9289 52742 9301 52794
rect 9353 52742 9365 52794
rect 9417 52742 10856 52794
rect 1104 52720 10856 52742
rect 3786 52680 3792 52692
rect 3747 52652 3792 52680
rect 3786 52640 3792 52652
rect 3844 52640 3850 52692
rect 290 52572 296 52624
rect 348 52612 354 52624
rect 1210 52612 1216 52624
rect 348 52584 1216 52612
rect 348 52572 354 52584
rect 1210 52572 1216 52584
rect 1268 52612 1274 52624
rect 2590 52612 2596 52624
rect 1268 52584 2596 52612
rect 1268 52572 1274 52584
rect 2590 52572 2596 52584
rect 2648 52572 2654 52624
rect 2777 52615 2835 52621
rect 2777 52581 2789 52615
rect 2823 52612 2835 52615
rect 2866 52612 2872 52624
rect 2823 52584 2872 52612
rect 2823 52581 2835 52584
rect 2777 52575 2835 52581
rect 2866 52572 2872 52584
rect 2924 52612 2930 52624
rect 3878 52612 3884 52624
rect 2924 52584 3884 52612
rect 2924 52572 2930 52584
rect 3878 52572 3884 52584
rect 3936 52612 3942 52624
rect 5166 52612 5172 52624
rect 3936 52584 5172 52612
rect 3936 52572 3942 52584
rect 5166 52572 5172 52584
rect 5224 52572 5230 52624
rect 9950 52544 9956 52556
rect 1780 52516 9956 52544
rect 842 52436 848 52488
rect 900 52436 906 52488
rect 1486 52436 1492 52488
rect 1544 52476 1550 52488
rect 1780 52485 1808 52516
rect 9950 52504 9956 52516
rect 10008 52504 10014 52556
rect 1581 52479 1639 52485
rect 1581 52476 1593 52479
rect 1544 52448 1593 52476
rect 1544 52436 1550 52448
rect 1581 52445 1593 52448
rect 1627 52445 1639 52479
rect 1581 52439 1639 52445
rect 1765 52479 1823 52485
rect 1765 52445 1777 52479
rect 1811 52445 1823 52479
rect 1946 52476 1952 52488
rect 1907 52448 1952 52476
rect 1765 52439 1823 52445
rect 1946 52436 1952 52448
rect 2004 52436 2010 52488
rect 2590 52476 2596 52488
rect 2551 52448 2596 52476
rect 2590 52436 2596 52448
rect 2648 52436 2654 52488
rect 3326 52436 3332 52488
rect 3384 52476 3390 52488
rect 3789 52479 3847 52485
rect 3789 52476 3801 52479
rect 3384 52448 3801 52476
rect 3384 52436 3390 52448
rect 3789 52445 3801 52448
rect 3835 52445 3847 52479
rect 3789 52439 3847 52445
rect 3973 52479 4031 52485
rect 3973 52445 3985 52479
rect 4019 52476 4031 52479
rect 4614 52476 4620 52488
rect 4019 52448 4620 52476
rect 4019 52445 4031 52448
rect 3973 52439 4031 52445
rect 4614 52436 4620 52448
rect 4672 52436 4678 52488
rect 860 52408 888 52436
rect 1673 52411 1731 52417
rect 860 52380 1532 52408
rect 845 52343 903 52349
rect 845 52309 857 52343
rect 891 52340 903 52343
rect 1397 52343 1455 52349
rect 1397 52340 1409 52343
rect 891 52312 1409 52340
rect 891 52309 903 52312
rect 845 52303 903 52309
rect 1397 52309 1409 52312
rect 1443 52309 1455 52343
rect 1504 52340 1532 52380
rect 1673 52377 1685 52411
rect 1719 52377 1731 52411
rect 1673 52371 1731 52377
rect 1688 52340 1716 52371
rect 2130 52368 2136 52420
rect 2188 52408 2194 52420
rect 2314 52408 2320 52420
rect 2188 52380 2320 52408
rect 2188 52368 2194 52380
rect 2314 52368 2320 52380
rect 2372 52368 2378 52420
rect 1504 52312 1716 52340
rect 1397 52303 1455 52309
rect 1104 52250 10856 52272
rect 1104 52198 4213 52250
rect 4265 52198 4277 52250
rect 4329 52198 4341 52250
rect 4393 52198 4405 52250
rect 4457 52198 4469 52250
rect 4521 52198 7477 52250
rect 7529 52198 7541 52250
rect 7593 52198 7605 52250
rect 7657 52198 7669 52250
rect 7721 52198 7733 52250
rect 7785 52198 10856 52250
rect 1104 52176 10856 52198
rect 937 52139 995 52145
rect 937 52105 949 52139
rect 983 52136 995 52139
rect 2130 52136 2136 52148
rect 983 52108 2136 52136
rect 983 52105 995 52108
rect 937 52099 995 52105
rect 2130 52096 2136 52108
rect 2188 52096 2194 52148
rect 2406 51960 2412 52012
rect 2464 52000 2470 52012
rect 2501 52003 2559 52009
rect 2501 52000 2513 52003
rect 2464 51972 2513 52000
rect 2464 51960 2470 51972
rect 2501 51969 2513 51972
rect 2547 51969 2559 52003
rect 10134 52000 10140 52012
rect 10095 51972 10140 52000
rect 2501 51963 2559 51969
rect 10134 51960 10140 51972
rect 10192 51960 10198 52012
rect 1486 51892 1492 51944
rect 1544 51932 1550 51944
rect 1854 51932 1860 51944
rect 1544 51904 1860 51932
rect 1544 51892 1550 51904
rect 1854 51892 1860 51904
rect 1912 51932 1918 51944
rect 2225 51935 2283 51941
rect 2225 51932 2237 51935
rect 1912 51904 2237 51932
rect 1912 51892 1918 51904
rect 2225 51901 2237 51904
rect 2271 51901 2283 51935
rect 2225 51895 2283 51901
rect 2961 51935 3019 51941
rect 2961 51901 2973 51935
rect 3007 51901 3019 51935
rect 2961 51895 3019 51901
rect 3237 51935 3295 51941
rect 3237 51901 3249 51935
rect 3283 51932 3295 51935
rect 3326 51932 3332 51944
rect 3283 51904 3332 51932
rect 3283 51901 3295 51904
rect 3237 51895 3295 51901
rect 2976 51864 3004 51895
rect 3326 51892 3332 51904
rect 3384 51892 3390 51944
rect 3694 51864 3700 51876
rect 2976 51836 3700 51864
rect 3694 51824 3700 51836
rect 3752 51864 3758 51876
rect 6638 51864 6644 51876
rect 3752 51836 6644 51864
rect 3752 51824 3758 51836
rect 6638 51824 6644 51836
rect 6696 51824 6702 51876
rect 937 51799 995 51805
rect 937 51765 949 51799
rect 983 51796 995 51799
rect 1578 51796 1584 51808
rect 983 51768 1584 51796
rect 983 51765 995 51768
rect 937 51759 995 51765
rect 1578 51756 1584 51768
rect 1636 51756 1642 51808
rect 9950 51796 9956 51808
rect 9911 51768 9956 51796
rect 9950 51756 9956 51768
rect 10008 51756 10014 51808
rect 1104 51706 10856 51728
rect 1104 51654 2582 51706
rect 2634 51654 2646 51706
rect 2698 51654 2710 51706
rect 2762 51654 2774 51706
rect 2826 51654 2838 51706
rect 2890 51654 5845 51706
rect 5897 51654 5909 51706
rect 5961 51654 5973 51706
rect 6025 51654 6037 51706
rect 6089 51654 6101 51706
rect 6153 51654 9109 51706
rect 9161 51654 9173 51706
rect 9225 51654 9237 51706
rect 9289 51654 9301 51706
rect 9353 51654 9365 51706
rect 9417 51654 10856 51706
rect 1104 51632 10856 51654
rect 1946 51592 1952 51604
rect 1504 51564 1952 51592
rect 1397 51391 1455 51397
rect 1397 51357 1409 51391
rect 1443 51388 1455 51391
rect 1504 51388 1532 51564
rect 1946 51552 1952 51564
rect 2004 51552 2010 51604
rect 3786 51552 3792 51604
rect 3844 51592 3850 51604
rect 9858 51592 9864 51604
rect 3844 51564 9864 51592
rect 3844 51552 3850 51564
rect 9858 51552 9864 51564
rect 9916 51552 9922 51604
rect 1964 51524 1992 51552
rect 1964 51496 2820 51524
rect 1443 51360 1532 51388
rect 1443 51357 1455 51360
rect 1397 51351 1455 51357
rect 1578 51348 1584 51400
rect 1636 51388 1642 51400
rect 1636 51360 1681 51388
rect 1636 51348 1642 51360
rect 1762 51348 1768 51400
rect 1820 51388 1826 51400
rect 2593 51391 2651 51397
rect 2593 51388 2605 51391
rect 1820 51360 2605 51388
rect 1820 51348 1826 51360
rect 2593 51357 2605 51360
rect 2639 51357 2651 51391
rect 2792 51388 2820 51496
rect 3694 51484 3700 51536
rect 3752 51524 3758 51536
rect 3970 51524 3976 51536
rect 3752 51496 3976 51524
rect 3752 51484 3758 51496
rect 3970 51484 3976 51496
rect 4028 51484 4034 51536
rect 5534 51484 5540 51536
rect 5592 51524 5598 51536
rect 5810 51524 5816 51536
rect 5592 51496 5816 51524
rect 5592 51484 5598 51496
rect 5810 51484 5816 51496
rect 5868 51484 5874 51536
rect 2961 51391 3019 51397
rect 2961 51388 2973 51391
rect 2792 51360 2973 51388
rect 2593 51351 2651 51357
rect 2961 51357 2973 51360
rect 3007 51357 3019 51391
rect 3786 51388 3792 51400
rect 3747 51360 3792 51388
rect 2961 51351 3019 51357
rect 3786 51348 3792 51360
rect 3844 51348 3850 51400
rect 1670 51320 1676 51332
rect 1631 51292 1676 51320
rect 1670 51280 1676 51292
rect 1728 51280 1734 51332
rect 2314 51280 2320 51332
rect 2372 51320 2378 51332
rect 2685 51323 2743 51329
rect 2685 51320 2697 51323
rect 2372 51292 2697 51320
rect 2372 51280 2378 51292
rect 2685 51289 2697 51292
rect 2731 51289 2743 51323
rect 2685 51283 2743 51289
rect 2777 51323 2835 51329
rect 2777 51289 2789 51323
rect 2823 51320 2835 51323
rect 9950 51320 9956 51332
rect 2823 51292 9956 51320
rect 2823 51289 2835 51292
rect 2777 51283 2835 51289
rect 9950 51280 9956 51292
rect 10008 51280 10014 51332
rect 1949 51255 2007 51261
rect 1949 51221 1961 51255
rect 1995 51252 2007 51255
rect 2130 51252 2136 51264
rect 1995 51224 2136 51252
rect 1995 51221 2007 51224
rect 1949 51215 2007 51221
rect 2130 51212 2136 51224
rect 2188 51212 2194 51264
rect 2409 51255 2467 51261
rect 2409 51221 2421 51255
rect 2455 51252 2467 51255
rect 2590 51252 2596 51264
rect 2455 51224 2596 51252
rect 2455 51221 2467 51224
rect 2409 51215 2467 51221
rect 2590 51212 2596 51224
rect 2648 51212 2654 51264
rect 3970 51252 3976 51264
rect 3931 51224 3976 51252
rect 3970 51212 3976 51224
rect 4028 51212 4034 51264
rect 1104 51162 10856 51184
rect 1104 51110 4213 51162
rect 4265 51110 4277 51162
rect 4329 51110 4341 51162
rect 4393 51110 4405 51162
rect 4457 51110 4469 51162
rect 4521 51110 7477 51162
rect 7529 51110 7541 51162
rect 7593 51110 7605 51162
rect 7657 51110 7669 51162
rect 7721 51110 7733 51162
rect 7785 51110 10856 51162
rect 1104 51088 10856 51110
rect 845 51051 903 51057
rect 845 51017 857 51051
rect 891 51048 903 51051
rect 1302 51048 1308 51060
rect 891 51020 1308 51048
rect 891 51017 903 51020
rect 845 51011 903 51017
rect 1302 51008 1308 51020
rect 1360 51008 1366 51060
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 3476 51020 3521 51048
rect 3476 51008 3482 51020
rect 9858 51008 9864 51060
rect 9916 51048 9922 51060
rect 9953 51051 10011 51057
rect 9953 51048 9965 51051
rect 9916 51020 9965 51048
rect 9916 51008 9922 51020
rect 9953 51017 9965 51020
rect 9999 51017 10011 51051
rect 9953 51011 10011 51017
rect 1949 50915 2007 50921
rect 1949 50881 1961 50915
rect 1995 50912 2007 50915
rect 2958 50912 2964 50924
rect 1995 50884 2964 50912
rect 1995 50881 2007 50884
rect 1949 50875 2007 50881
rect 2958 50872 2964 50884
rect 3016 50872 3022 50924
rect 3262 50915 3320 50921
rect 3262 50881 3274 50915
rect 3308 50912 3320 50915
rect 3973 50915 4031 50921
rect 3308 50884 3832 50912
rect 3308 50881 3320 50884
rect 3262 50875 3320 50881
rect 1854 50804 1860 50856
rect 1912 50844 1918 50856
rect 2225 50847 2283 50853
rect 2225 50844 2237 50847
rect 1912 50816 2237 50844
rect 1912 50804 1918 50816
rect 2225 50813 2237 50816
rect 2271 50813 2283 50847
rect 2225 50807 2283 50813
rect 1670 50736 1676 50788
rect 1728 50776 1734 50788
rect 2590 50776 2596 50788
rect 1728 50748 2596 50776
rect 1728 50736 1734 50748
rect 2590 50736 2596 50748
rect 2648 50736 2654 50788
rect 3050 50736 3056 50788
rect 3108 50776 3114 50788
rect 3804 50776 3832 50884
rect 3973 50881 3985 50915
rect 4019 50881 4031 50915
rect 3973 50875 4031 50881
rect 4157 50915 4215 50921
rect 4157 50881 4169 50915
rect 4203 50912 4215 50915
rect 5166 50912 5172 50924
rect 4203 50884 5172 50912
rect 4203 50881 4215 50884
rect 4157 50875 4215 50881
rect 3878 50804 3884 50856
rect 3936 50844 3942 50856
rect 3988 50844 4016 50875
rect 5166 50872 5172 50884
rect 5224 50872 5230 50924
rect 5534 50872 5540 50924
rect 5592 50872 5598 50924
rect 10134 50912 10140 50924
rect 10095 50884 10140 50912
rect 10134 50872 10140 50884
rect 10192 50872 10198 50924
rect 3936 50816 4016 50844
rect 3936 50804 3942 50816
rect 4154 50776 4160 50788
rect 3108 50748 3464 50776
rect 3804 50748 4160 50776
rect 3108 50736 3114 50748
rect 3436 50708 3464 50748
rect 4154 50736 4160 50748
rect 4212 50736 4218 50788
rect 3973 50711 4031 50717
rect 3973 50708 3985 50711
rect 3436 50680 3985 50708
rect 3973 50677 3985 50680
rect 4019 50677 4031 50711
rect 3973 50671 4031 50677
rect 5442 50668 5448 50720
rect 5500 50708 5506 50720
rect 5552 50708 5580 50872
rect 5810 50736 5816 50788
rect 5868 50776 5874 50788
rect 6730 50776 6736 50788
rect 5868 50748 6736 50776
rect 5868 50736 5874 50748
rect 6730 50736 6736 50748
rect 6788 50736 6794 50788
rect 5500 50680 5580 50708
rect 5500 50668 5506 50680
rect 1104 50618 10856 50640
rect 1104 50566 2582 50618
rect 2634 50566 2646 50618
rect 2698 50566 2710 50618
rect 2762 50566 2774 50618
rect 2826 50566 2838 50618
rect 2890 50566 5845 50618
rect 5897 50566 5909 50618
rect 5961 50566 5973 50618
rect 6025 50566 6037 50618
rect 6089 50566 6101 50618
rect 6153 50566 9109 50618
rect 9161 50566 9173 50618
rect 9225 50566 9237 50618
rect 9289 50566 9301 50618
rect 9353 50566 9365 50618
rect 9417 50566 10856 50618
rect 1104 50544 10856 50566
rect 1762 50368 1768 50380
rect 1596 50340 1768 50368
rect 1596 50309 1624 50340
rect 1762 50328 1768 50340
rect 1820 50328 1826 50380
rect 3326 50328 3332 50380
rect 3384 50368 3390 50380
rect 3786 50368 3792 50380
rect 3384 50340 3792 50368
rect 3384 50328 3390 50340
rect 3786 50328 3792 50340
rect 3844 50328 3850 50380
rect 3878 50328 3884 50380
rect 3936 50368 3942 50380
rect 4065 50371 4123 50377
rect 4065 50368 4077 50371
rect 3936 50340 4077 50368
rect 3936 50328 3942 50340
rect 4065 50337 4077 50340
rect 4111 50337 4123 50371
rect 4065 50331 4123 50337
rect 1581 50303 1639 50309
rect 1581 50269 1593 50303
rect 1627 50269 1639 50303
rect 1581 50263 1639 50269
rect 1854 50260 1860 50312
rect 1912 50300 1918 50312
rect 1949 50303 2007 50309
rect 1949 50300 1961 50303
rect 1912 50272 1961 50300
rect 1912 50260 1918 50272
rect 1949 50269 1961 50272
rect 1995 50269 2007 50303
rect 1949 50263 2007 50269
rect 2590 50260 2596 50312
rect 2648 50300 2654 50312
rect 2685 50303 2743 50309
rect 2685 50300 2697 50303
rect 2648 50272 2697 50300
rect 2648 50260 2654 50272
rect 2685 50269 2697 50272
rect 2731 50269 2743 50303
rect 2685 50263 2743 50269
rect 3234 50260 3240 50312
rect 3292 50300 3298 50312
rect 4154 50300 4160 50312
rect 3292 50272 4160 50300
rect 3292 50260 3298 50272
rect 4154 50260 4160 50272
rect 4212 50260 4218 50312
rect 1673 50235 1731 50241
rect 1673 50201 1685 50235
rect 1719 50201 1731 50235
rect 1673 50195 1731 50201
rect 1765 50235 1823 50241
rect 1765 50201 1777 50235
rect 1811 50232 1823 50235
rect 9950 50232 9956 50244
rect 1811 50204 9956 50232
rect 1811 50201 1823 50204
rect 1765 50195 1823 50201
rect 1210 50124 1216 50176
rect 1268 50164 1274 50176
rect 1397 50167 1455 50173
rect 1397 50164 1409 50167
rect 1268 50136 1409 50164
rect 1268 50124 1274 50136
rect 1397 50133 1409 50136
rect 1443 50133 1455 50167
rect 1688 50164 1716 50195
rect 9950 50192 9956 50204
rect 10008 50192 10014 50244
rect 1946 50164 1952 50176
rect 1688 50136 1952 50164
rect 1397 50127 1455 50133
rect 1946 50124 1952 50136
rect 2004 50124 2010 50176
rect 2498 50164 2504 50176
rect 2459 50136 2504 50164
rect 2498 50124 2504 50136
rect 2556 50124 2562 50176
rect 1104 50074 10856 50096
rect 1104 50022 4213 50074
rect 4265 50022 4277 50074
rect 4329 50022 4341 50074
rect 4393 50022 4405 50074
rect 4457 50022 4469 50074
rect 4521 50022 7477 50074
rect 7529 50022 7541 50074
rect 7593 50022 7605 50074
rect 7657 50022 7669 50074
rect 7721 50022 7733 50074
rect 7785 50022 10856 50074
rect 1104 50000 10856 50022
rect 1486 49960 1492 49972
rect 1447 49932 1492 49960
rect 1486 49920 1492 49932
rect 1544 49920 1550 49972
rect 2961 49963 3019 49969
rect 1688 49932 2774 49960
rect 1688 49833 1716 49932
rect 2746 49892 2774 49932
rect 2961 49929 2973 49963
rect 3007 49960 3019 49963
rect 3694 49960 3700 49972
rect 3007 49932 3700 49960
rect 3007 49929 3019 49932
rect 2961 49923 3019 49929
rect 3694 49920 3700 49932
rect 3752 49920 3758 49972
rect 9950 49960 9956 49972
rect 9911 49932 9956 49960
rect 9950 49920 9956 49932
rect 10008 49920 10014 49972
rect 3605 49895 3663 49901
rect 3605 49892 3617 49895
rect 2746 49864 3617 49892
rect 3605 49861 3617 49864
rect 3651 49861 3663 49895
rect 3605 49855 3663 49861
rect 1673 49827 1731 49833
rect 1673 49793 1685 49827
rect 1719 49793 1731 49827
rect 1673 49787 1731 49793
rect 2409 49827 2467 49833
rect 2409 49793 2421 49827
rect 2455 49824 2467 49827
rect 2455 49796 2636 49824
rect 2455 49793 2467 49796
rect 2409 49787 2467 49793
rect 1946 49716 1952 49768
rect 2004 49756 2010 49768
rect 2222 49756 2228 49768
rect 2004 49728 2228 49756
rect 2004 49716 2010 49728
rect 2222 49716 2228 49728
rect 2280 49716 2286 49768
rect 2608 49756 2636 49796
rect 2682 49784 2688 49836
rect 2740 49824 2746 49836
rect 2869 49827 2927 49833
rect 2869 49824 2881 49827
rect 2740 49796 2881 49824
rect 2740 49784 2746 49796
rect 2869 49793 2881 49796
rect 2915 49793 2927 49827
rect 2869 49787 2927 49793
rect 2958 49784 2964 49836
rect 3016 49824 3022 49836
rect 3053 49827 3111 49833
rect 3053 49824 3065 49827
rect 3016 49796 3065 49824
rect 3016 49784 3022 49796
rect 3053 49793 3065 49796
rect 3099 49824 3111 49827
rect 3513 49827 3571 49833
rect 3513 49824 3525 49827
rect 3099 49796 3525 49824
rect 3099 49793 3111 49796
rect 3053 49787 3111 49793
rect 3513 49793 3525 49796
rect 3559 49793 3571 49827
rect 3513 49787 3571 49793
rect 3697 49827 3755 49833
rect 3697 49793 3709 49827
rect 3743 49824 3755 49827
rect 6454 49824 6460 49836
rect 3743 49796 6460 49824
rect 3743 49793 3755 49796
rect 3697 49787 3755 49793
rect 3418 49756 3424 49768
rect 2608 49728 3424 49756
rect 3418 49716 3424 49728
rect 3476 49716 3482 49768
rect 3528 49756 3556 49787
rect 6454 49784 6460 49796
rect 6512 49784 6518 49836
rect 10137 49827 10195 49833
rect 10137 49793 10149 49827
rect 10183 49793 10195 49827
rect 10137 49787 10195 49793
rect 3878 49756 3884 49768
rect 3528 49728 3884 49756
rect 3878 49716 3884 49728
rect 3936 49716 3942 49768
rect 10152 49700 10180 49787
rect 198 49648 204 49700
rect 256 49688 262 49700
rect 2682 49688 2688 49700
rect 256 49660 2688 49688
rect 256 49648 262 49660
rect 2682 49648 2688 49660
rect 2740 49648 2746 49700
rect 2866 49648 2872 49700
rect 2924 49688 2930 49700
rect 3694 49688 3700 49700
rect 2924 49660 3700 49688
rect 2924 49648 2930 49660
rect 3694 49648 3700 49660
rect 3752 49648 3758 49700
rect 10134 49648 10140 49700
rect 10192 49648 10198 49700
rect 2222 49620 2228 49632
rect 2183 49592 2228 49620
rect 2222 49580 2228 49592
rect 2280 49580 2286 49632
rect 1104 49530 10856 49552
rect 1104 49478 2582 49530
rect 2634 49478 2646 49530
rect 2698 49478 2710 49530
rect 2762 49478 2774 49530
rect 2826 49478 2838 49530
rect 2890 49478 5845 49530
rect 5897 49478 5909 49530
rect 5961 49478 5973 49530
rect 6025 49478 6037 49530
rect 6089 49478 6101 49530
rect 6153 49478 9109 49530
rect 9161 49478 9173 49530
rect 9225 49478 9237 49530
rect 9289 49478 9301 49530
rect 9353 49478 9365 49530
rect 9417 49478 10856 49530
rect 1104 49456 10856 49478
rect 1394 49376 1400 49428
rect 1452 49416 1458 49428
rect 1854 49416 1860 49428
rect 1452 49388 1860 49416
rect 1452 49376 1458 49388
rect 1854 49376 1860 49388
rect 1912 49376 1918 49428
rect 2593 49419 2651 49425
rect 2593 49385 2605 49419
rect 2639 49416 2651 49419
rect 3234 49416 3240 49428
rect 2639 49388 3240 49416
rect 2639 49385 2651 49388
rect 2593 49379 2651 49385
rect 3234 49376 3240 49388
rect 3292 49376 3298 49428
rect 753 49351 811 49357
rect 753 49317 765 49351
rect 799 49348 811 49351
rect 3053 49351 3111 49357
rect 3053 49348 3065 49351
rect 799 49320 3065 49348
rect 799 49317 811 49320
rect 753 49311 811 49317
rect 3053 49317 3065 49320
rect 3099 49317 3111 49351
rect 3053 49311 3111 49317
rect 1118 49240 1124 49292
rect 1176 49280 1182 49292
rect 1394 49280 1400 49292
rect 1176 49252 1400 49280
rect 1176 49240 1182 49252
rect 1394 49240 1400 49252
rect 1452 49240 1458 49292
rect 2774 49280 2780 49292
rect 2424 49252 2780 49280
rect 2424 49221 2452 49252
rect 2774 49240 2780 49252
rect 2832 49240 2838 49292
rect 3786 49280 3792 49292
rect 3747 49252 3792 49280
rect 3786 49240 3792 49252
rect 3844 49240 3850 49292
rect 1673 49215 1731 49221
rect 1673 49181 1685 49215
rect 1719 49181 1731 49215
rect 1673 49175 1731 49181
rect 2409 49215 2467 49221
rect 2409 49181 2421 49215
rect 2455 49181 2467 49215
rect 2409 49175 2467 49181
rect 2593 49215 2651 49221
rect 2593 49181 2605 49215
rect 2639 49212 2651 49215
rect 2958 49212 2964 49224
rect 2639 49184 2964 49212
rect 2639 49181 2651 49184
rect 2593 49175 2651 49181
rect 1118 49104 1124 49156
rect 1176 49144 1182 49156
rect 1688 49144 1716 49175
rect 2958 49172 2964 49184
rect 3016 49212 3022 49224
rect 3053 49215 3111 49221
rect 3053 49212 3065 49215
rect 3016 49184 3065 49212
rect 3016 49172 3022 49184
rect 3053 49181 3065 49184
rect 3099 49181 3111 49215
rect 3053 49175 3111 49181
rect 3237 49215 3295 49221
rect 3237 49181 3249 49215
rect 3283 49181 3295 49215
rect 3237 49175 3295 49181
rect 2866 49144 2872 49156
rect 1176 49116 1624 49144
rect 1688 49116 2872 49144
rect 1176 49104 1182 49116
rect 1486 49076 1492 49088
rect 1447 49048 1492 49076
rect 1486 49036 1492 49048
rect 1544 49036 1550 49088
rect 1596 49076 1624 49116
rect 2866 49104 2872 49116
rect 2924 49104 2930 49156
rect 3252 49144 3280 49175
rect 3878 49172 3884 49224
rect 3936 49212 3942 49224
rect 4065 49215 4123 49221
rect 4065 49212 4077 49215
rect 3936 49184 4077 49212
rect 3936 49172 3942 49184
rect 4065 49181 4077 49184
rect 4111 49181 4123 49215
rect 4065 49175 4123 49181
rect 2976 49116 3280 49144
rect 2976 49076 3004 49116
rect 1596 49048 3004 49076
rect 1104 48986 10856 49008
rect 1104 48934 4213 48986
rect 4265 48934 4277 48986
rect 4329 48934 4341 48986
rect 4393 48934 4405 48986
rect 4457 48934 4469 48986
rect 4521 48934 7477 48986
rect 7529 48934 7541 48986
rect 7593 48934 7605 48986
rect 7657 48934 7669 48986
rect 7721 48934 7733 48986
rect 7785 48934 10856 48986
rect 1104 48912 10856 48934
rect 2774 48764 2780 48816
rect 2832 48804 2838 48816
rect 4522 48804 4528 48816
rect 2832 48776 4528 48804
rect 2832 48764 2838 48776
rect 4522 48764 4528 48776
rect 4580 48764 4586 48816
rect 1673 48739 1731 48745
rect 1673 48705 1685 48739
rect 1719 48705 1731 48739
rect 1673 48699 1731 48705
rect 2409 48739 2467 48745
rect 2409 48705 2421 48739
rect 2455 48736 2467 48739
rect 3694 48736 3700 48748
rect 2455 48708 3700 48736
rect 2455 48705 2467 48708
rect 2409 48699 2467 48705
rect 1688 48668 1716 48699
rect 3694 48696 3700 48708
rect 3752 48696 3758 48748
rect 10134 48736 10140 48748
rect 10095 48708 10140 48736
rect 10134 48696 10140 48708
rect 10192 48696 10198 48748
rect 6822 48668 6828 48680
rect 1688 48640 6828 48668
rect 6822 48628 6828 48640
rect 6880 48628 6886 48680
rect 2222 48600 2228 48612
rect 2183 48572 2228 48600
rect 2222 48560 2228 48572
rect 2280 48560 2286 48612
rect 1486 48532 1492 48544
rect 1447 48504 1492 48532
rect 1486 48492 1492 48504
rect 1544 48492 1550 48544
rect 9953 48535 10011 48541
rect 9953 48501 9965 48535
rect 9999 48532 10011 48535
rect 10965 48535 11023 48541
rect 10965 48532 10977 48535
rect 9999 48504 10977 48532
rect 9999 48501 10011 48504
rect 9953 48495 10011 48501
rect 10965 48501 10977 48504
rect 11011 48501 11023 48535
rect 10965 48495 11023 48501
rect 1104 48442 10856 48464
rect 1104 48390 2582 48442
rect 2634 48390 2646 48442
rect 2698 48390 2710 48442
rect 2762 48390 2774 48442
rect 2826 48390 2838 48442
rect 2890 48390 5845 48442
rect 5897 48390 5909 48442
rect 5961 48390 5973 48442
rect 6025 48390 6037 48442
rect 6089 48390 6101 48442
rect 6153 48390 9109 48442
rect 9161 48390 9173 48442
rect 9225 48390 9237 48442
rect 9289 48390 9301 48442
rect 9353 48390 9365 48442
rect 9417 48390 10856 48442
rect 1104 48368 10856 48390
rect 937 48331 995 48337
rect 937 48297 949 48331
rect 983 48328 995 48331
rect 1762 48328 1768 48340
rect 983 48300 1768 48328
rect 983 48297 995 48300
rect 937 48291 995 48297
rect 1762 48288 1768 48300
rect 1820 48288 1826 48340
rect 2498 48260 2504 48272
rect 2459 48232 2504 48260
rect 2498 48220 2504 48232
rect 2556 48220 2562 48272
rect 750 48152 756 48204
rect 808 48192 814 48204
rect 808 48164 2728 48192
rect 808 48152 814 48164
rect 1670 48124 1676 48136
rect 1631 48096 1676 48124
rect 1670 48084 1676 48096
rect 1728 48084 1734 48136
rect 2700 48133 2728 48164
rect 2501 48127 2559 48133
rect 2501 48093 2513 48127
rect 2547 48093 2559 48127
rect 2501 48087 2559 48093
rect 2685 48127 2743 48133
rect 2685 48093 2697 48127
rect 2731 48093 2743 48127
rect 2685 48087 2743 48093
rect 2516 48056 2544 48087
rect 2866 48056 2872 48068
rect 2516 48028 2872 48056
rect 2866 48016 2872 48028
rect 2924 48016 2930 48068
rect 1486 47988 1492 48000
rect 1447 47960 1492 47988
rect 1486 47948 1492 47960
rect 1544 47948 1550 48000
rect 2774 47948 2780 48000
rect 2832 47988 2838 48000
rect 3326 47988 3332 48000
rect 2832 47960 3332 47988
rect 2832 47948 2838 47960
rect 3326 47948 3332 47960
rect 3384 47948 3390 48000
rect 1104 47898 10856 47920
rect 1104 47846 4213 47898
rect 4265 47846 4277 47898
rect 4329 47846 4341 47898
rect 4393 47846 4405 47898
rect 4457 47846 4469 47898
rect 4521 47846 7477 47898
rect 7529 47846 7541 47898
rect 7593 47846 7605 47898
rect 7657 47846 7669 47898
rect 7721 47846 7733 47898
rect 7785 47846 10856 47898
rect 1104 47824 10856 47846
rect 658 47744 664 47796
rect 716 47784 722 47796
rect 3326 47784 3332 47796
rect 716 47756 3332 47784
rect 716 47744 722 47756
rect 3326 47744 3332 47756
rect 3384 47744 3390 47796
rect 2958 47676 2964 47728
rect 3016 47716 3022 47728
rect 3016 47688 3061 47716
rect 3016 47676 3022 47688
rect 1394 47608 1400 47660
rect 1452 47648 1458 47660
rect 1673 47651 1731 47657
rect 1673 47648 1685 47651
rect 1452 47620 1685 47648
rect 1452 47608 1458 47620
rect 1673 47617 1685 47620
rect 1719 47617 1731 47651
rect 1673 47611 1731 47617
rect 2409 47651 2467 47657
rect 2409 47617 2421 47651
rect 2455 47648 2467 47651
rect 2774 47648 2780 47660
rect 2455 47620 2780 47648
rect 2455 47617 2467 47620
rect 2409 47611 2467 47617
rect 2774 47608 2780 47620
rect 2832 47608 2838 47660
rect 2866 47608 2872 47660
rect 2924 47648 2930 47660
rect 3053 47651 3111 47657
rect 2924 47620 2969 47648
rect 2924 47608 2930 47620
rect 3053 47617 3065 47651
rect 3099 47617 3111 47651
rect 10134 47648 10140 47660
rect 10095 47620 10140 47648
rect 3053 47611 3111 47617
rect 842 47472 848 47524
rect 900 47512 906 47524
rect 3068 47512 3096 47611
rect 10134 47608 10140 47620
rect 10192 47608 10198 47660
rect 900 47484 3096 47512
rect 900 47472 906 47484
rect 1486 47444 1492 47456
rect 1447 47416 1492 47444
rect 1486 47404 1492 47416
rect 1544 47404 1550 47456
rect 2222 47444 2228 47456
rect 2183 47416 2228 47444
rect 2222 47404 2228 47416
rect 2280 47404 2286 47456
rect 9953 47447 10011 47453
rect 9953 47413 9965 47447
rect 9999 47444 10011 47447
rect 11057 47447 11115 47453
rect 11057 47444 11069 47447
rect 9999 47416 11069 47444
rect 9999 47413 10011 47416
rect 9953 47407 10011 47413
rect 11057 47413 11069 47416
rect 11103 47413 11115 47447
rect 11057 47407 11115 47413
rect 1104 47354 10856 47376
rect 1104 47302 2582 47354
rect 2634 47302 2646 47354
rect 2698 47302 2710 47354
rect 2762 47302 2774 47354
rect 2826 47302 2838 47354
rect 2890 47302 5845 47354
rect 5897 47302 5909 47354
rect 5961 47302 5973 47354
rect 6025 47302 6037 47354
rect 6089 47302 6101 47354
rect 6153 47302 9109 47354
rect 9161 47302 9173 47354
rect 9225 47302 9237 47354
rect 9289 47302 9301 47354
rect 9353 47302 9365 47354
rect 9417 47302 10856 47354
rect 1104 47280 10856 47302
rect 1670 47200 1676 47252
rect 1728 47240 1734 47252
rect 2501 47243 2559 47249
rect 2501 47240 2513 47243
rect 1728 47212 2513 47240
rect 1728 47200 1734 47212
rect 2501 47209 2513 47212
rect 2547 47209 2559 47243
rect 2501 47203 2559 47209
rect 3418 47200 3424 47252
rect 3476 47240 3482 47252
rect 3789 47243 3847 47249
rect 3789 47240 3801 47243
rect 3476 47212 3801 47240
rect 3476 47200 3482 47212
rect 3789 47209 3801 47212
rect 3835 47209 3847 47243
rect 3789 47203 3847 47209
rect 4890 47172 4896 47184
rect 1688 47144 4896 47172
rect 1026 47064 1032 47116
rect 1084 47064 1090 47116
rect 1044 47036 1072 47064
rect 1578 47036 1584 47048
rect 1044 47008 1584 47036
rect 1578 46996 1584 47008
rect 1636 46996 1642 47048
rect 1688 47045 1716 47144
rect 4890 47132 4896 47144
rect 4948 47132 4954 47184
rect 2516 47076 3832 47104
rect 2516 47045 2544 47076
rect 3804 47045 3832 47076
rect 1673 47039 1731 47045
rect 1673 47005 1685 47039
rect 1719 47005 1731 47039
rect 1673 46999 1731 47005
rect 2501 47039 2559 47045
rect 2501 47005 2513 47039
rect 2547 47005 2559 47039
rect 2501 46999 2559 47005
rect 2685 47039 2743 47045
rect 2685 47005 2697 47039
rect 2731 47005 2743 47039
rect 2685 46999 2743 47005
rect 3789 47039 3847 47045
rect 3789 47005 3801 47039
rect 3835 47036 3847 47039
rect 3878 47036 3884 47048
rect 3835 47008 3884 47036
rect 3835 47005 3847 47008
rect 3789 46999 3847 47005
rect 2700 46968 2728 46999
rect 3878 46996 3884 47008
rect 3936 46996 3942 47048
rect 3973 47039 4031 47045
rect 3973 47005 3985 47039
rect 4019 47005 4031 47039
rect 3973 46999 4031 47005
rect 1044 46940 2728 46968
rect 198 46764 204 46776
rect 159 46736 204 46764
rect 198 46724 204 46736
rect 256 46724 262 46776
rect 1044 46696 1072 46940
rect 2958 46928 2964 46980
rect 3016 46968 3022 46980
rect 3988 46968 4016 46999
rect 3016 46940 4016 46968
rect 3016 46928 3022 46940
rect 1302 46860 1308 46912
rect 1360 46900 1366 46912
rect 1489 46903 1547 46909
rect 1489 46900 1501 46903
rect 1360 46872 1501 46900
rect 1360 46860 1366 46872
rect 1489 46869 1501 46872
rect 1535 46869 1547 46903
rect 1489 46863 1547 46869
rect 2774 46860 2780 46912
rect 2832 46900 2838 46912
rect 8294 46900 8300 46912
rect 2832 46872 8300 46900
rect 2832 46860 2838 46872
rect 8294 46860 8300 46872
rect 8352 46860 8358 46912
rect 1104 46810 10856 46832
rect 1104 46758 4213 46810
rect 4265 46758 4277 46810
rect 4329 46758 4341 46810
rect 4393 46758 4405 46810
rect 4457 46758 4469 46810
rect 4521 46758 7477 46810
rect 7529 46758 7541 46810
rect 7593 46758 7605 46810
rect 7657 46758 7669 46810
rect 7721 46758 7733 46810
rect 7785 46758 10856 46810
rect 1104 46736 10856 46758
rect 1118 46696 1124 46708
rect 1044 46668 1124 46696
rect 1118 46656 1124 46668
rect 1176 46656 1182 46708
rect 3694 46696 3700 46708
rect 3655 46668 3700 46696
rect 3694 46656 3700 46668
rect 3752 46656 3758 46708
rect 198 46588 204 46640
rect 256 46628 262 46640
rect 3878 46628 3884 46640
rect 256 46600 1808 46628
rect 256 46588 262 46600
rect 1673 46563 1731 46569
rect 1673 46529 1685 46563
rect 1719 46529 1731 46563
rect 1673 46523 1731 46529
rect 1688 46424 1716 46523
rect 1780 46492 1808 46600
rect 3620 46600 3884 46628
rect 2409 46563 2467 46569
rect 2409 46529 2421 46563
rect 2455 46560 2467 46563
rect 2774 46560 2780 46572
rect 2455 46532 2780 46560
rect 2455 46529 2467 46532
rect 2409 46523 2467 46529
rect 2774 46520 2780 46532
rect 2832 46520 2838 46572
rect 2869 46563 2927 46569
rect 2869 46529 2881 46563
rect 2915 46560 2927 46563
rect 3050 46560 3056 46572
rect 2915 46532 3056 46560
rect 2915 46529 2927 46532
rect 2869 46523 2927 46529
rect 3050 46520 3056 46532
rect 3108 46520 3114 46572
rect 3620 46569 3648 46600
rect 3878 46588 3884 46600
rect 3936 46588 3942 46640
rect 3605 46563 3663 46569
rect 3605 46529 3617 46563
rect 3651 46529 3663 46563
rect 3605 46523 3663 46529
rect 3789 46563 3847 46569
rect 3789 46529 3801 46563
rect 3835 46529 3847 46563
rect 10134 46560 10140 46572
rect 10095 46532 10140 46560
rect 3789 46523 3847 46529
rect 3804 46492 3832 46523
rect 10134 46520 10140 46532
rect 10192 46520 10198 46572
rect 1780 46464 3832 46492
rect 3050 46424 3056 46436
rect 1688 46396 2774 46424
rect 3011 46396 3056 46424
rect 1394 46316 1400 46368
rect 1452 46356 1458 46368
rect 1489 46359 1547 46365
rect 1489 46356 1501 46359
rect 1452 46328 1501 46356
rect 1452 46316 1458 46328
rect 1489 46325 1501 46328
rect 1535 46325 1547 46359
rect 2222 46356 2228 46368
rect 2183 46328 2228 46356
rect 1489 46319 1547 46325
rect 2222 46316 2228 46328
rect 2280 46316 2286 46368
rect 2746 46356 2774 46396
rect 3050 46384 3056 46396
rect 3108 46384 3114 46436
rect 6730 46424 6736 46436
rect 3160 46396 6736 46424
rect 3160 46356 3188 46396
rect 6730 46384 6736 46396
rect 6788 46384 6794 46436
rect 2746 46328 3188 46356
rect 4614 46316 4620 46368
rect 4672 46356 4678 46368
rect 4890 46356 4896 46368
rect 4672 46328 4896 46356
rect 4672 46316 4678 46328
rect 4890 46316 4896 46328
rect 4948 46316 4954 46368
rect 9950 46356 9956 46368
rect 9911 46328 9956 46356
rect 9950 46316 9956 46328
rect 10008 46316 10014 46368
rect 1104 46266 10856 46288
rect 290 46180 296 46232
rect 348 46220 354 46232
rect 658 46220 664 46232
rect 348 46192 664 46220
rect 348 46180 354 46192
rect 658 46180 664 46192
rect 716 46180 722 46232
rect 1104 46214 2582 46266
rect 2634 46214 2646 46266
rect 2698 46214 2710 46266
rect 2762 46214 2774 46266
rect 2826 46214 2838 46266
rect 2890 46214 5845 46266
rect 5897 46214 5909 46266
rect 5961 46214 5973 46266
rect 6025 46214 6037 46266
rect 6089 46214 6101 46266
rect 6153 46214 9109 46266
rect 9161 46214 9173 46266
rect 9225 46214 9237 46266
rect 9289 46214 9301 46266
rect 9353 46214 9365 46266
rect 9417 46214 10856 46266
rect 1104 46192 10856 46214
rect 106 46112 112 46164
rect 164 46152 170 46164
rect 3050 46152 3056 46164
rect 164 46124 3056 46152
rect 164 46112 170 46124
rect 3050 46112 3056 46124
rect 3108 46112 3114 46164
rect 3234 46112 3240 46164
rect 3292 46112 3298 46164
rect 4614 46112 4620 46164
rect 4672 46152 4678 46164
rect 5074 46152 5080 46164
rect 4672 46124 5080 46152
rect 4672 46112 4678 46124
rect 5074 46112 5080 46124
rect 5132 46112 5138 46164
rect 201 46087 259 46093
rect 201 46053 213 46087
rect 247 46084 259 46087
rect 290 46084 296 46096
rect 247 46056 296 46084
rect 247 46053 259 46056
rect 201 46047 259 46053
rect 290 46044 296 46056
rect 348 46044 354 46096
rect 2406 46016 2412 46028
rect 2367 45988 2412 46016
rect 2406 45976 2412 45988
rect 2464 45976 2470 46028
rect 3252 46016 3280 46112
rect 3160 45988 3280 46016
rect 3160 45960 3188 45988
rect 3326 45976 3332 46028
rect 3384 46016 3390 46028
rect 3510 46016 3516 46028
rect 3384 45988 3516 46016
rect 3384 45976 3390 45988
rect 3510 45976 3516 45988
rect 3568 45976 3574 46028
rect 1578 45908 1584 45960
rect 1636 45948 1642 45960
rect 1673 45951 1731 45957
rect 1673 45948 1685 45951
rect 1636 45920 1685 45948
rect 1636 45908 1642 45920
rect 1673 45917 1685 45920
rect 1719 45917 1731 45951
rect 1673 45911 1731 45917
rect 2685 45951 2743 45957
rect 2685 45917 2697 45951
rect 2731 45917 2743 45951
rect 2685 45911 2743 45917
rect 1486 45812 1492 45824
rect 1447 45784 1492 45812
rect 1486 45772 1492 45784
rect 1544 45772 1550 45824
rect 2222 45772 2228 45824
rect 2280 45812 2286 45824
rect 2700 45812 2728 45911
rect 3142 45908 3148 45960
rect 3200 45908 3206 45960
rect 3234 45908 3240 45960
rect 3292 45948 3298 45960
rect 3694 45948 3700 45960
rect 3292 45920 3700 45948
rect 3292 45908 3298 45920
rect 3694 45908 3700 45920
rect 3752 45908 3758 45960
rect 2280 45784 2728 45812
rect 2280 45772 2286 45784
rect 1104 45722 10856 45744
rect 1104 45670 4213 45722
rect 4265 45670 4277 45722
rect 4329 45670 4341 45722
rect 4393 45670 4405 45722
rect 4457 45670 4469 45722
rect 4521 45670 7477 45722
rect 7529 45670 7541 45722
rect 7593 45670 7605 45722
rect 7657 45670 7669 45722
rect 7721 45670 7733 45722
rect 7785 45670 10856 45722
rect 1104 45648 10856 45670
rect 382 45568 388 45620
rect 440 45608 446 45620
rect 1578 45608 1584 45620
rect 440 45580 1584 45608
rect 440 45568 446 45580
rect 1578 45568 1584 45580
rect 1636 45568 1642 45620
rect 3326 45500 3332 45552
rect 3384 45540 3390 45552
rect 5534 45540 5540 45552
rect 3384 45512 5540 45540
rect 3384 45500 3390 45512
rect 5534 45500 5540 45512
rect 5592 45500 5598 45552
rect 2685 45475 2743 45481
rect 2685 45441 2697 45475
rect 2731 45472 2743 45475
rect 3970 45472 3976 45484
rect 2731 45444 3976 45472
rect 2731 45441 2743 45444
rect 2685 45435 2743 45441
rect 3970 45432 3976 45444
rect 4028 45432 4034 45484
rect 10134 45472 10140 45484
rect 10095 45444 10140 45472
rect 10134 45432 10140 45444
rect 10192 45432 10198 45484
rect 2406 45404 2412 45416
rect 2367 45376 2412 45404
rect 2406 45364 2412 45376
rect 2464 45364 2470 45416
rect 9858 45228 9864 45280
rect 9916 45268 9922 45280
rect 9953 45271 10011 45277
rect 9953 45268 9965 45271
rect 9916 45240 9965 45268
rect 9916 45228 9922 45240
rect 9953 45237 9965 45240
rect 9999 45237 10011 45271
rect 9953 45231 10011 45237
rect 1104 45178 10856 45200
rect 1104 45126 2582 45178
rect 2634 45126 2646 45178
rect 2698 45126 2710 45178
rect 2762 45126 2774 45178
rect 2826 45126 2838 45178
rect 2890 45126 5845 45178
rect 5897 45126 5909 45178
rect 5961 45126 5973 45178
rect 6025 45126 6037 45178
rect 6089 45126 6101 45178
rect 6153 45126 9109 45178
rect 9161 45126 9173 45178
rect 9225 45126 9237 45178
rect 9289 45126 9301 45178
rect 9353 45126 9365 45178
rect 9417 45126 10856 45178
rect 1104 45104 10856 45126
rect 1302 45024 1308 45076
rect 1360 45064 1366 45076
rect 2958 45064 2964 45076
rect 1360 45036 2964 45064
rect 1360 45024 1366 45036
rect 2958 45024 2964 45036
rect 3016 45024 3022 45076
rect 2222 44928 2228 44940
rect 1596 44900 2228 44928
rect 1596 44869 1624 44900
rect 2222 44888 2228 44900
rect 2280 44928 2286 44940
rect 2590 44928 2596 44940
rect 2280 44900 2596 44928
rect 2280 44888 2286 44900
rect 2590 44888 2596 44900
rect 2648 44888 2654 44940
rect 1581 44863 1639 44869
rect 1581 44829 1593 44863
rect 1627 44829 1639 44863
rect 1581 44823 1639 44829
rect 1949 44863 2007 44869
rect 1949 44829 1961 44863
rect 1995 44860 2007 44863
rect 2406 44860 2412 44872
rect 1995 44832 2412 44860
rect 1995 44829 2007 44832
rect 1949 44823 2007 44829
rect 2406 44820 2412 44832
rect 2464 44820 2470 44872
rect 2685 44863 2743 44869
rect 2685 44829 2697 44863
rect 2731 44860 2743 44863
rect 3786 44860 3792 44872
rect 2731 44832 3792 44860
rect 2731 44829 2743 44832
rect 2685 44823 2743 44829
rect 3786 44820 3792 44832
rect 3844 44820 3850 44872
rect 937 44795 995 44801
rect 937 44761 949 44795
rect 983 44792 995 44795
rect 1673 44795 1731 44801
rect 1673 44792 1685 44795
rect 983 44764 1685 44792
rect 983 44761 995 44764
rect 937 44755 995 44761
rect 1673 44761 1685 44764
rect 1719 44761 1731 44795
rect 1673 44755 1731 44761
rect 1765 44795 1823 44801
rect 1765 44761 1777 44795
rect 1811 44792 1823 44795
rect 11057 44795 11115 44801
rect 11057 44792 11069 44795
rect 1811 44764 11069 44792
rect 1811 44761 1823 44764
rect 1765 44755 1823 44761
rect 11057 44761 11069 44764
rect 11103 44761 11115 44795
rect 11057 44755 11115 44761
rect 1394 44724 1400 44736
rect 1355 44696 1400 44724
rect 1394 44684 1400 44696
rect 1452 44684 1458 44736
rect 1578 44684 1584 44736
rect 1636 44724 1642 44736
rect 2501 44727 2559 44733
rect 2501 44724 2513 44727
rect 1636 44696 2513 44724
rect 1636 44684 1642 44696
rect 2501 44693 2513 44696
rect 2547 44693 2559 44727
rect 2501 44687 2559 44693
rect 1104 44634 10856 44656
rect 1104 44582 4213 44634
rect 4265 44582 4277 44634
rect 4329 44582 4341 44634
rect 4393 44582 4405 44634
rect 4457 44582 4469 44634
rect 4521 44582 7477 44634
rect 7529 44582 7541 44634
rect 7593 44582 7605 44634
rect 7657 44582 7669 44634
rect 7721 44582 7733 44634
rect 7785 44582 10856 44634
rect 1104 44560 10856 44582
rect 2590 44520 2596 44532
rect 1504 44492 2596 44520
rect 106 44412 112 44464
rect 164 44452 170 44464
rect 842 44452 848 44464
rect 164 44424 848 44452
rect 164 44412 170 44424
rect 842 44412 848 44424
rect 900 44412 906 44464
rect 1504 44396 1532 44492
rect 2590 44480 2596 44492
rect 2648 44480 2654 44532
rect 10965 44523 11023 44529
rect 10965 44520 10977 44523
rect 2792 44492 10977 44520
rect 1670 44452 1676 44464
rect 1631 44424 1676 44452
rect 1670 44412 1676 44424
rect 1728 44412 1734 44464
rect 2498 44412 2504 44464
rect 2556 44452 2562 44464
rect 2792 44461 2820 44492
rect 10965 44489 10977 44492
rect 11011 44489 11023 44523
rect 10965 44483 11023 44489
rect 2685 44455 2743 44461
rect 2685 44452 2697 44455
rect 2556 44424 2697 44452
rect 2556 44412 2562 44424
rect 2685 44421 2697 44424
rect 2731 44421 2743 44455
rect 2685 44415 2743 44421
rect 2777 44455 2835 44461
rect 2777 44421 2789 44455
rect 2823 44421 2835 44455
rect 9950 44452 9956 44464
rect 2777 44415 2835 44421
rect 2884 44424 9956 44452
rect 1486 44384 1492 44396
rect 1399 44356 1492 44384
rect 1486 44344 1492 44356
rect 1544 44384 1550 44396
rect 1581 44387 1639 44393
rect 1581 44384 1593 44387
rect 1544 44356 1593 44384
rect 1544 44344 1550 44356
rect 1581 44353 1593 44356
rect 1627 44353 1639 44387
rect 1581 44347 1639 44353
rect 1765 44387 1823 44393
rect 1765 44353 1777 44387
rect 1811 44353 1823 44387
rect 1765 44347 1823 44353
rect 1949 44387 2007 44393
rect 1949 44353 1961 44387
rect 1995 44384 2007 44387
rect 2406 44384 2412 44396
rect 1995 44356 2412 44384
rect 1995 44353 2007 44356
rect 1949 44347 2007 44353
rect 1780 44316 1808 44347
rect 2406 44344 2412 44356
rect 2464 44344 2470 44396
rect 2590 44384 2596 44396
rect 2551 44356 2596 44384
rect 2590 44344 2596 44356
rect 2648 44344 2654 44396
rect 2884 44316 2912 44424
rect 9950 44412 9956 44424
rect 10008 44412 10014 44464
rect 2961 44387 3019 44393
rect 2961 44353 2973 44387
rect 3007 44384 3019 44387
rect 10134 44384 10140 44396
rect 3007 44356 3096 44384
rect 10095 44356 10140 44384
rect 3007 44353 3019 44356
rect 2961 44347 3019 44353
rect 1780 44288 2912 44316
rect 2498 44208 2504 44260
rect 2556 44248 2562 44260
rect 3068 44248 3096 44356
rect 10134 44344 10140 44356
rect 10192 44344 10198 44396
rect 2556 44220 3096 44248
rect 2556 44208 2562 44220
rect 1397 44183 1455 44189
rect 1397 44149 1409 44183
rect 1443 44180 1455 44183
rect 1854 44180 1860 44192
rect 1443 44152 1860 44180
rect 1443 44149 1455 44152
rect 1397 44143 1455 44149
rect 1854 44140 1860 44152
rect 1912 44140 1918 44192
rect 2406 44180 2412 44192
rect 2367 44152 2412 44180
rect 2406 44140 2412 44152
rect 2464 44140 2470 44192
rect 9950 44180 9956 44192
rect 9911 44152 9956 44180
rect 9950 44140 9956 44152
rect 10008 44140 10014 44192
rect 1104 44090 10856 44112
rect 1104 44038 2582 44090
rect 2634 44038 2646 44090
rect 2698 44038 2710 44090
rect 2762 44038 2774 44090
rect 2826 44038 2838 44090
rect 2890 44038 5845 44090
rect 5897 44038 5909 44090
rect 5961 44038 5973 44090
rect 6025 44038 6037 44090
rect 6089 44038 6101 44090
rect 6153 44038 9109 44090
rect 9161 44038 9173 44090
rect 9225 44038 9237 44090
rect 9289 44038 9301 44090
rect 9353 44038 9365 44090
rect 9417 44038 10856 44090
rect 1104 44016 10856 44038
rect 2498 43840 2504 43852
rect 1964 43812 2504 43840
rect 1486 43732 1492 43784
rect 1544 43772 1550 43784
rect 1581 43775 1639 43781
rect 1581 43772 1593 43775
rect 1544 43744 1593 43772
rect 1544 43732 1550 43744
rect 1581 43741 1593 43744
rect 1627 43741 1639 43775
rect 1581 43735 1639 43741
rect 1670 43732 1676 43784
rect 1728 43772 1734 43784
rect 1964 43781 1992 43812
rect 2498 43800 2504 43812
rect 2556 43800 2562 43852
rect 1949 43775 2007 43781
rect 1728 43744 1773 43772
rect 1728 43732 1734 43744
rect 1949 43741 1961 43775
rect 1995 43741 2007 43775
rect 1949 43735 2007 43741
rect 2222 43732 2228 43784
rect 2280 43772 2286 43784
rect 2409 43775 2467 43781
rect 2409 43772 2421 43775
rect 2280 43744 2421 43772
rect 2280 43732 2286 43744
rect 2409 43741 2421 43744
rect 2455 43741 2467 43775
rect 2409 43735 2467 43741
rect 3789 43775 3847 43781
rect 3789 43741 3801 43775
rect 3835 43772 3847 43775
rect 4062 43772 4068 43784
rect 3835 43744 4068 43772
rect 3835 43741 3847 43744
rect 3789 43735 3847 43741
rect 4062 43732 4068 43744
rect 4120 43732 4126 43784
rect 1765 43707 1823 43713
rect 1765 43673 1777 43707
rect 1811 43704 1823 43707
rect 9950 43704 9956 43716
rect 1811 43676 9956 43704
rect 1811 43673 1823 43676
rect 1765 43667 1823 43673
rect 9950 43664 9956 43676
rect 10008 43664 10014 43716
rect 1397 43639 1455 43645
rect 1397 43605 1409 43639
rect 1443 43636 1455 43639
rect 1578 43636 1584 43648
rect 1443 43608 1584 43636
rect 1443 43605 1455 43608
rect 1397 43599 1455 43605
rect 1578 43596 1584 43608
rect 1636 43596 1642 43648
rect 2593 43639 2651 43645
rect 2593 43605 2605 43639
rect 2639 43636 2651 43639
rect 2774 43636 2780 43648
rect 2639 43608 2780 43636
rect 2639 43605 2651 43608
rect 2593 43599 2651 43605
rect 2774 43596 2780 43608
rect 2832 43596 2838 43648
rect 3970 43636 3976 43648
rect 3931 43608 3976 43636
rect 3970 43596 3976 43608
rect 4028 43596 4034 43648
rect 1104 43546 10856 43568
rect 1104 43494 4213 43546
rect 4265 43494 4277 43546
rect 4329 43494 4341 43546
rect 4393 43494 4405 43546
rect 4457 43494 4469 43546
rect 4521 43494 7477 43546
rect 7529 43494 7541 43546
rect 7593 43494 7605 43546
rect 7657 43494 7669 43546
rect 7721 43494 7733 43546
rect 7785 43494 10856 43546
rect 1104 43472 10856 43494
rect 9858 43432 9864 43444
rect 1780 43404 9864 43432
rect 1780 43373 1808 43404
rect 9858 43392 9864 43404
rect 9916 43392 9922 43444
rect 1765 43367 1823 43373
rect 1765 43333 1777 43367
rect 1811 43333 1823 43367
rect 1765 43327 1823 43333
rect 4154 43324 4160 43376
rect 4212 43364 4218 43376
rect 4982 43364 4988 43376
rect 4212 43336 4988 43364
rect 4212 43324 4218 43336
rect 4982 43324 4988 43336
rect 5040 43324 5046 43376
rect 1486 43256 1492 43308
rect 1544 43296 1550 43308
rect 1581 43299 1639 43305
rect 1581 43296 1593 43299
rect 1544 43268 1593 43296
rect 1544 43256 1550 43268
rect 1581 43265 1593 43268
rect 1627 43265 1639 43299
rect 1581 43259 1639 43265
rect 1673 43299 1731 43305
rect 1673 43265 1685 43299
rect 1719 43265 1731 43299
rect 1673 43259 1731 43265
rect 1949 43299 2007 43305
rect 1949 43265 1961 43299
rect 1995 43296 2007 43299
rect 2498 43296 2504 43308
rect 1995 43268 2504 43296
rect 1995 43265 2007 43268
rect 1949 43259 2007 43265
rect 1688 43228 1716 43259
rect 2498 43256 2504 43268
rect 2556 43256 2562 43308
rect 2685 43299 2743 43305
rect 2685 43265 2697 43299
rect 2731 43296 2743 43299
rect 3142 43296 3148 43308
rect 2731 43268 3148 43296
rect 2731 43265 2743 43268
rect 2685 43259 2743 43265
rect 3142 43256 3148 43268
rect 3200 43256 3206 43308
rect 9858 43296 9864 43308
rect 9819 43268 9864 43296
rect 9858 43256 9864 43268
rect 9916 43256 9922 43308
rect 8478 43228 8484 43240
rect 1688 43200 8484 43228
rect 8478 43188 8484 43200
rect 8536 43188 8542 43240
rect 937 43095 995 43101
rect 937 43061 949 43095
rect 983 43092 995 43095
rect 1397 43095 1455 43101
rect 1397 43092 1409 43095
rect 983 43064 1409 43092
rect 983 43061 995 43064
rect 937 43055 995 43061
rect 1397 43061 1409 43064
rect 1443 43061 1455 43095
rect 2498 43092 2504 43104
rect 2459 43064 2504 43092
rect 1397 43055 1455 43061
rect 2498 43052 2504 43064
rect 2556 43052 2562 43104
rect 10042 43092 10048 43104
rect 10003 43064 10048 43092
rect 10042 43052 10048 43064
rect 10100 43052 10106 43104
rect 1104 43002 10856 43024
rect 1104 42950 2582 43002
rect 2634 42950 2646 43002
rect 2698 42950 2710 43002
rect 2762 42950 2774 43002
rect 2826 42950 2838 43002
rect 2890 42950 5845 43002
rect 5897 42950 5909 43002
rect 5961 42950 5973 43002
rect 6025 42950 6037 43002
rect 6089 42950 6101 43002
rect 6153 42950 9109 43002
rect 9161 42950 9173 43002
rect 9225 42950 9237 43002
rect 9289 42950 9301 43002
rect 9353 42950 9365 43002
rect 9417 42950 10856 43002
rect 1104 42928 10856 42950
rect 4709 42891 4767 42897
rect 4709 42857 4721 42891
rect 4755 42888 4767 42891
rect 4755 42860 5304 42888
rect 4755 42857 4767 42860
rect 4709 42851 4767 42857
rect 14 42780 20 42832
rect 72 42820 78 42832
rect 72 42792 1072 42820
rect 72 42780 78 42792
rect 934 42712 940 42764
rect 992 42712 998 42764
rect 14 42644 20 42696
rect 72 42684 78 42696
rect 750 42684 756 42696
rect 72 42656 756 42684
rect 72 42644 78 42656
rect 750 42644 756 42656
rect 808 42644 814 42696
rect 952 42492 980 42712
rect 934 42440 940 42492
rect 992 42440 998 42492
rect 290 42372 296 42424
rect 348 42412 354 42424
rect 842 42412 848 42424
rect 348 42384 848 42412
rect 348 42372 354 42384
rect 842 42372 848 42384
rect 900 42372 906 42424
rect 1044 42344 1072 42792
rect 5276 42752 5304 42860
rect 9858 42752 9864 42764
rect 2746 42724 5120 42752
rect 5276 42724 9864 42752
rect 1670 42684 1676 42696
rect 1631 42656 1676 42684
rect 1670 42644 1676 42656
rect 1728 42644 1734 42696
rect 2409 42687 2467 42693
rect 2409 42653 2421 42687
rect 2455 42684 2467 42687
rect 2746 42684 2774 42724
rect 2455 42656 2774 42684
rect 4525 42687 4583 42693
rect 2455 42653 2467 42656
rect 2409 42647 2467 42653
rect 4525 42653 4537 42687
rect 4571 42653 4583 42687
rect 4525 42647 4583 42653
rect 4709 42687 4767 42693
rect 4709 42653 4721 42687
rect 4755 42684 4767 42687
rect 4982 42684 4988 42696
rect 4755 42656 4988 42684
rect 4755 42653 4767 42656
rect 4709 42647 4767 42653
rect 4540 42616 4568 42647
rect 4982 42644 4988 42656
rect 5040 42644 5046 42696
rect 5092 42684 5120 42724
rect 9858 42712 9864 42724
rect 9916 42712 9922 42764
rect 8386 42684 8392 42696
rect 5092 42656 8392 42684
rect 8386 42644 8392 42656
rect 8444 42644 8450 42696
rect 5442 42616 5448 42628
rect 4540 42588 5448 42616
rect 5442 42576 5448 42588
rect 5500 42576 5506 42628
rect 1486 42548 1492 42560
rect 1447 42520 1492 42548
rect 1486 42508 1492 42520
rect 1544 42508 1550 42560
rect 2222 42548 2228 42560
rect 2183 42520 2228 42548
rect 2222 42508 2228 42520
rect 2280 42508 2286 42560
rect 1104 42458 10856 42480
rect 1104 42406 4213 42458
rect 4265 42406 4277 42458
rect 4329 42406 4341 42458
rect 4393 42406 4405 42458
rect 4457 42406 4469 42458
rect 4521 42406 7477 42458
rect 7529 42406 7541 42458
rect 7593 42406 7605 42458
rect 7657 42406 7669 42458
rect 7721 42406 7733 42458
rect 7785 42406 10856 42458
rect 1104 42384 10856 42406
rect 1044 42316 1440 42344
rect 845 42279 903 42285
rect 845 42245 857 42279
rect 891 42276 903 42279
rect 1412 42276 1440 42316
rect 1670 42304 1676 42356
rect 1728 42344 1734 42356
rect 6914 42344 6920 42356
rect 1728 42316 6920 42344
rect 1728 42304 1734 42316
rect 6914 42304 6920 42316
rect 6972 42304 6978 42356
rect 4890 42276 4896 42288
rect 891 42248 980 42276
rect 1412 42248 1716 42276
rect 891 42245 903 42248
rect 845 42239 903 42245
rect 952 42208 980 42248
rect 1688 42217 1716 42248
rect 4540 42248 4896 42276
rect 4540 42217 4568 42248
rect 4890 42236 4896 42248
rect 4948 42276 4954 42288
rect 5074 42276 5080 42288
rect 4948 42248 5080 42276
rect 4948 42236 4954 42248
rect 5074 42236 5080 42248
rect 5132 42236 5138 42288
rect 1673 42211 1731 42217
rect 952 42180 1624 42208
rect 1596 42152 1624 42180
rect 1673 42177 1685 42211
rect 1719 42177 1731 42211
rect 1673 42171 1731 42177
rect 4525 42211 4583 42217
rect 4525 42177 4537 42211
rect 4571 42177 4583 42211
rect 4525 42171 4583 42177
rect 4709 42211 4767 42217
rect 4709 42177 4721 42211
rect 4755 42208 4767 42211
rect 4982 42208 4988 42220
rect 4755 42180 4988 42208
rect 4755 42177 4767 42180
rect 4709 42171 4767 42177
rect 4982 42168 4988 42180
rect 5040 42168 5046 42220
rect 9861 42211 9919 42217
rect 9861 42177 9873 42211
rect 9907 42177 9919 42211
rect 9861 42171 9919 42177
rect 845 42143 903 42149
rect 845 42109 857 42143
rect 891 42140 903 42143
rect 1394 42140 1400 42152
rect 891 42112 1400 42140
rect 891 42109 903 42112
rect 845 42103 903 42109
rect 1394 42100 1400 42112
rect 1452 42100 1458 42152
rect 1578 42100 1584 42152
rect 1636 42100 1642 42152
rect 4617 42143 4675 42149
rect 4617 42109 4629 42143
rect 4663 42140 4675 42143
rect 9876 42140 9904 42171
rect 4663 42112 9904 42140
rect 4663 42109 4675 42112
rect 4617 42103 4675 42109
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 1489 42007 1547 42013
rect 1489 42004 1501 42007
rect 1452 41976 1501 42004
rect 1452 41964 1458 41976
rect 1489 41973 1501 41976
rect 1535 41973 1547 42007
rect 10042 42004 10048 42016
rect 10003 41976 10048 42004
rect 1489 41967 1547 41973
rect 10042 41964 10048 41976
rect 10100 41964 10106 42016
rect 1104 41914 10856 41936
rect 1104 41862 2582 41914
rect 2634 41862 2646 41914
rect 2698 41862 2710 41914
rect 2762 41862 2774 41914
rect 2826 41862 2838 41914
rect 2890 41862 5845 41914
rect 5897 41862 5909 41914
rect 5961 41862 5973 41914
rect 6025 41862 6037 41914
rect 6089 41862 6101 41914
rect 6153 41862 9109 41914
rect 9161 41862 9173 41914
rect 9225 41862 9237 41914
rect 9289 41862 9301 41914
rect 9353 41862 9365 41914
rect 9417 41862 10856 41914
rect 1104 41840 10856 41862
rect 1946 41692 1952 41744
rect 2004 41732 2010 41744
rect 2314 41732 2320 41744
rect 2004 41704 2320 41732
rect 2004 41692 2010 41704
rect 2314 41692 2320 41704
rect 2372 41692 2378 41744
rect 1673 41599 1731 41605
rect 1673 41565 1685 41599
rect 1719 41596 1731 41599
rect 6730 41596 6736 41608
rect 1719 41568 6736 41596
rect 1719 41565 1731 41568
rect 1673 41559 1731 41565
rect 6730 41556 6736 41568
rect 6788 41556 6794 41608
rect 1210 41488 1216 41540
rect 1268 41528 1274 41540
rect 1946 41528 1952 41540
rect 1268 41500 1952 41528
rect 1268 41488 1274 41500
rect 1946 41488 1952 41500
rect 2004 41488 2010 41540
rect 3786 41488 3792 41540
rect 3844 41528 3850 41540
rect 5258 41528 5264 41540
rect 3844 41500 5264 41528
rect 3844 41488 3850 41500
rect 5258 41488 5264 41500
rect 5316 41488 5322 41540
rect 1486 41460 1492 41472
rect 1447 41432 1492 41460
rect 1486 41420 1492 41432
rect 1544 41420 1550 41472
rect 1104 41370 10856 41392
rect 1104 41318 4213 41370
rect 4265 41318 4277 41370
rect 4329 41318 4341 41370
rect 4393 41318 4405 41370
rect 4457 41318 4469 41370
rect 4521 41318 7477 41370
rect 7529 41318 7541 41370
rect 7593 41318 7605 41370
rect 7657 41318 7669 41370
rect 7721 41318 7733 41370
rect 7785 41318 10856 41370
rect 1104 41296 10856 41318
rect 8570 41256 8576 41268
rect 1688 41228 8576 41256
rect 1688 41129 1716 41228
rect 8570 41216 8576 41228
rect 8628 41216 8634 41268
rect 4890 41188 4896 41200
rect 4540 41160 4896 41188
rect 4540 41129 4568 41160
rect 4890 41148 4896 41160
rect 4948 41188 4954 41200
rect 5350 41188 5356 41200
rect 4948 41160 5356 41188
rect 4948 41148 4954 41160
rect 5350 41148 5356 41160
rect 5408 41148 5414 41200
rect 1673 41123 1731 41129
rect 1673 41089 1685 41123
rect 1719 41089 1731 41123
rect 1673 41083 1731 41089
rect 4525 41123 4583 41129
rect 4525 41089 4537 41123
rect 4571 41089 4583 41123
rect 4525 41083 4583 41089
rect 4709 41123 4767 41129
rect 4709 41089 4721 41123
rect 4755 41120 4767 41123
rect 4982 41120 4988 41132
rect 4755 41092 4988 41120
rect 4755 41089 4767 41092
rect 4709 41083 4767 41089
rect 4982 41080 4988 41092
rect 5040 41080 5046 41132
rect 9861 41123 9919 41129
rect 9861 41120 9873 41123
rect 6886 41092 9873 41120
rect 1486 40916 1492 40928
rect 1447 40888 1492 40916
rect 1486 40876 1492 40888
rect 1544 40876 1550 40928
rect 4709 40919 4767 40925
rect 4709 40885 4721 40919
rect 4755 40916 4767 40919
rect 6886 40916 6914 41092
rect 9861 41089 9873 41092
rect 9907 41089 9919 41123
rect 9861 41083 9919 41089
rect 10042 40916 10048 40928
rect 4755 40888 6914 40916
rect 10003 40888 10048 40916
rect 4755 40885 4767 40888
rect 4709 40879 4767 40885
rect 10042 40876 10048 40888
rect 10100 40876 10106 40928
rect 1104 40826 10856 40848
rect 1104 40774 2582 40826
rect 2634 40774 2646 40826
rect 2698 40774 2710 40826
rect 2762 40774 2774 40826
rect 2826 40774 2838 40826
rect 2890 40774 5845 40826
rect 5897 40774 5909 40826
rect 5961 40774 5973 40826
rect 6025 40774 6037 40826
rect 6089 40774 6101 40826
rect 6153 40774 9109 40826
rect 9161 40774 9173 40826
rect 9225 40774 9237 40826
rect 9289 40774 9301 40826
rect 9353 40774 9365 40826
rect 9417 40774 10856 40826
rect 1104 40752 10856 40774
rect 106 40672 112 40724
rect 164 40712 170 40724
rect 1302 40712 1308 40724
rect 164 40684 1308 40712
rect 164 40672 170 40684
rect 1302 40672 1308 40684
rect 1360 40672 1366 40724
rect 3418 40672 3424 40724
rect 3476 40712 3482 40724
rect 3970 40712 3976 40724
rect 3476 40684 3976 40712
rect 3476 40672 3482 40684
rect 3970 40672 3976 40684
rect 4028 40672 4034 40724
rect 4798 40672 4804 40724
rect 4856 40712 4862 40724
rect 5350 40712 5356 40724
rect 4856 40684 5356 40712
rect 4856 40672 4862 40684
rect 5350 40672 5356 40684
rect 5408 40672 5414 40724
rect 290 40604 296 40656
rect 348 40644 354 40656
rect 1118 40644 1124 40656
rect 348 40616 1124 40644
rect 348 40604 354 40616
rect 1118 40604 1124 40616
rect 1176 40604 1182 40656
rect 1026 40536 1032 40588
rect 1084 40576 1090 40588
rect 1394 40576 1400 40588
rect 1084 40548 1400 40576
rect 1084 40536 1090 40548
rect 1394 40536 1400 40548
rect 1452 40536 1458 40588
rect 1673 40511 1731 40517
rect 1673 40477 1685 40511
rect 1719 40508 1731 40511
rect 8662 40508 8668 40520
rect 1719 40480 8668 40508
rect 1719 40477 1731 40480
rect 1673 40471 1731 40477
rect 8662 40468 8668 40480
rect 8720 40468 8726 40520
rect 1394 40400 1400 40452
rect 1452 40440 1458 40452
rect 2498 40440 2504 40452
rect 1452 40412 2504 40440
rect 1452 40400 1458 40412
rect 2498 40400 2504 40412
rect 2556 40400 2562 40452
rect 1486 40372 1492 40384
rect 1447 40344 1492 40372
rect 1486 40332 1492 40344
rect 1544 40332 1550 40384
rect 2406 40332 2412 40384
rect 2464 40372 2470 40384
rect 3786 40372 3792 40384
rect 2464 40344 3792 40372
rect 2464 40332 2470 40344
rect 3786 40332 3792 40344
rect 3844 40332 3850 40384
rect 1104 40282 10856 40304
rect 1104 40230 4213 40282
rect 4265 40230 4277 40282
rect 4329 40230 4341 40282
rect 4393 40230 4405 40282
rect 4457 40230 4469 40282
rect 4521 40230 7477 40282
rect 7529 40230 7541 40282
rect 7593 40230 7605 40282
rect 7657 40230 7669 40282
rect 7721 40230 7733 40282
rect 7785 40230 10856 40282
rect 1104 40208 10856 40230
rect 1670 40128 1676 40180
rect 1728 40168 1734 40180
rect 1854 40168 1860 40180
rect 1728 40140 1860 40168
rect 1728 40128 1734 40140
rect 1854 40128 1860 40140
rect 1912 40128 1918 40180
rect 2593 40171 2651 40177
rect 2593 40137 2605 40171
rect 2639 40168 2651 40171
rect 4614 40168 4620 40180
rect 2639 40140 4620 40168
rect 2639 40137 2651 40140
rect 2593 40131 2651 40137
rect 4614 40128 4620 40140
rect 4672 40128 4678 40180
rect 2406 40100 2412 40112
rect 1688 40072 2412 40100
rect 1688 40041 1716 40072
rect 2406 40060 2412 40072
rect 2464 40060 2470 40112
rect 4798 40100 4804 40112
rect 2700 40072 4804 40100
rect 1673 40035 1731 40041
rect 1673 40001 1685 40035
rect 1719 40001 1731 40035
rect 2498 40032 2504 40044
rect 2459 40004 2504 40032
rect 1673 39995 1731 40001
rect 2498 39992 2504 40004
rect 2556 39992 2562 40044
rect 2700 40041 2728 40072
rect 4798 40060 4804 40072
rect 4856 40060 4862 40112
rect 2685 40035 2743 40041
rect 2685 40001 2697 40035
rect 2731 40001 2743 40035
rect 2685 39995 2743 40001
rect 1486 39828 1492 39840
rect 1447 39800 1492 39828
rect 1486 39788 1492 39800
rect 1544 39788 1550 39840
rect 1104 39738 10856 39760
rect 1104 39686 2582 39738
rect 2634 39686 2646 39738
rect 2698 39686 2710 39738
rect 2762 39686 2774 39738
rect 2826 39686 2838 39738
rect 2890 39686 5845 39738
rect 5897 39686 5909 39738
rect 5961 39686 5973 39738
rect 6025 39686 6037 39738
rect 6089 39686 6101 39738
rect 6153 39686 9109 39738
rect 9161 39686 9173 39738
rect 9225 39686 9237 39738
rect 9289 39686 9301 39738
rect 9353 39686 9365 39738
rect 9417 39686 10856 39738
rect 1104 39664 10856 39686
rect 2409 39559 2467 39565
rect 2409 39525 2421 39559
rect 2455 39556 2467 39559
rect 5718 39556 5724 39568
rect 2455 39528 5724 39556
rect 2455 39525 2467 39528
rect 2409 39519 2467 39525
rect 5718 39516 5724 39528
rect 5776 39516 5782 39568
rect 3234 39488 3240 39500
rect 1688 39460 3240 39488
rect 1688 39429 1716 39460
rect 3234 39448 3240 39460
rect 3292 39448 3298 39500
rect 1673 39423 1731 39429
rect 1673 39389 1685 39423
rect 1719 39389 1731 39423
rect 2498 39420 2504 39432
rect 2459 39392 2504 39420
rect 1673 39383 1731 39389
rect 2498 39380 2504 39392
rect 2556 39380 2562 39432
rect 2685 39423 2743 39429
rect 2685 39389 2697 39423
rect 2731 39420 2743 39423
rect 2958 39420 2964 39432
rect 2731 39392 2964 39420
rect 2731 39389 2743 39392
rect 2685 39383 2743 39389
rect 2958 39380 2964 39392
rect 3016 39380 3022 39432
rect 9858 39420 9864 39432
rect 9819 39392 9864 39420
rect 9858 39380 9864 39392
rect 9916 39380 9922 39432
rect 1486 39284 1492 39296
rect 1447 39256 1492 39284
rect 1486 39244 1492 39256
rect 1544 39244 1550 39296
rect 10042 39284 10048 39296
rect 10003 39256 10048 39284
rect 10042 39244 10048 39256
rect 10100 39244 10106 39296
rect 1104 39194 10856 39216
rect 1104 39142 4213 39194
rect 4265 39142 4277 39194
rect 4329 39142 4341 39194
rect 4393 39142 4405 39194
rect 4457 39142 4469 39194
rect 4521 39142 7477 39194
rect 7529 39142 7541 39194
rect 7593 39142 7605 39194
rect 7657 39142 7669 39194
rect 7721 39142 7733 39194
rect 7785 39142 10856 39194
rect 1104 39120 10856 39142
rect 934 38972 940 39024
rect 992 39012 998 39024
rect 2317 39015 2375 39021
rect 2317 39012 2329 39015
rect 992 38984 2329 39012
rect 992 38972 998 38984
rect 2317 38981 2329 38984
rect 2363 38981 2375 39015
rect 2317 38975 2375 38981
rect 2406 38972 2412 39024
rect 2464 39012 2470 39024
rect 2464 38984 2636 39012
rect 2464 38972 2470 38984
rect 1578 38904 1584 38956
rect 1636 38944 1642 38956
rect 1673 38947 1731 38953
rect 1673 38944 1685 38947
rect 1636 38916 1685 38944
rect 1636 38904 1642 38916
rect 1673 38913 1685 38916
rect 1719 38913 1731 38947
rect 2498 38944 2504 38956
rect 2459 38916 2504 38944
rect 1673 38907 1731 38913
rect 2498 38904 2504 38916
rect 2556 38904 2562 38956
rect 2608 38953 2636 38984
rect 2593 38947 2651 38953
rect 2593 38913 2605 38947
rect 2639 38913 2651 38947
rect 2593 38907 2651 38913
rect 4249 38947 4307 38953
rect 4249 38913 4261 38947
rect 4295 38913 4307 38947
rect 4249 38907 4307 38913
rect 4433 38947 4491 38953
rect 4433 38913 4445 38947
rect 4479 38944 4491 38947
rect 4614 38944 4620 38956
rect 4479 38916 4620 38944
rect 4479 38913 4491 38916
rect 4433 38907 4491 38913
rect 4264 38876 4292 38907
rect 4614 38904 4620 38916
rect 4672 38904 4678 38956
rect 4798 38876 4804 38888
rect 4264 38848 4804 38876
rect 4798 38836 4804 38848
rect 4856 38836 4862 38888
rect 1486 38808 1492 38820
rect 1447 38780 1492 38808
rect 1486 38768 1492 38780
rect 1544 38768 1550 38820
rect 2958 38700 2964 38752
rect 3016 38740 3022 38752
rect 4246 38740 4252 38752
rect 3016 38712 4252 38740
rect 3016 38700 3022 38712
rect 4246 38700 4252 38712
rect 4304 38700 4310 38752
rect 4433 38743 4491 38749
rect 4433 38709 4445 38743
rect 4479 38740 4491 38743
rect 9858 38740 9864 38752
rect 4479 38712 9864 38740
rect 4479 38709 4491 38712
rect 4433 38703 4491 38709
rect 9858 38700 9864 38712
rect 9916 38700 9922 38752
rect 1104 38650 10856 38672
rect 1104 38598 2582 38650
rect 2634 38598 2646 38650
rect 2698 38598 2710 38650
rect 2762 38598 2774 38650
rect 2826 38598 2838 38650
rect 2890 38598 5845 38650
rect 5897 38598 5909 38650
rect 5961 38598 5973 38650
rect 6025 38598 6037 38650
rect 6089 38598 6101 38650
rect 6153 38598 9109 38650
rect 9161 38598 9173 38650
rect 9225 38598 9237 38650
rect 9289 38598 9301 38650
rect 9353 38598 9365 38650
rect 9417 38598 10856 38650
rect 1104 38576 10856 38598
rect 2409 38471 2467 38477
rect 2409 38437 2421 38471
rect 2455 38468 2467 38471
rect 7374 38468 7380 38480
rect 2455 38440 7380 38468
rect 2455 38437 2467 38440
rect 2409 38431 2467 38437
rect 7374 38428 7380 38440
rect 7432 38428 7438 38480
rect 2222 38400 2228 38412
rect 1688 38372 2228 38400
rect 1688 38341 1716 38372
rect 2222 38360 2228 38372
rect 2280 38360 2286 38412
rect 1673 38335 1731 38341
rect 1673 38301 1685 38335
rect 1719 38301 1731 38335
rect 2498 38332 2504 38344
rect 2459 38304 2504 38332
rect 1673 38295 1731 38301
rect 2498 38292 2504 38304
rect 2556 38292 2562 38344
rect 2593 38335 2651 38341
rect 2593 38301 2605 38335
rect 2639 38301 2651 38335
rect 4246 38332 4252 38344
rect 4207 38304 4252 38332
rect 2593 38295 2651 38301
rect 2222 38224 2228 38276
rect 2280 38264 2286 38276
rect 2608 38264 2636 38295
rect 4246 38292 4252 38304
rect 4304 38292 4310 38344
rect 4433 38335 4491 38341
rect 4433 38301 4445 38335
rect 4479 38332 4491 38335
rect 4614 38332 4620 38344
rect 4479 38304 4620 38332
rect 4479 38301 4491 38304
rect 4433 38295 4491 38301
rect 4614 38292 4620 38304
rect 4672 38292 4678 38344
rect 9861 38335 9919 38341
rect 9861 38332 9873 38335
rect 6886 38304 9873 38332
rect 2280 38236 2636 38264
rect 2280 38224 2286 38236
rect 1486 38196 1492 38208
rect 1447 38168 1492 38196
rect 1486 38156 1492 38168
rect 1544 38156 1550 38208
rect 4341 38199 4399 38205
rect 4341 38165 4353 38199
rect 4387 38196 4399 38199
rect 6886 38196 6914 38304
rect 9861 38301 9873 38304
rect 9907 38301 9919 38335
rect 9861 38295 9919 38301
rect 10042 38196 10048 38208
rect 4387 38168 6914 38196
rect 10003 38168 10048 38196
rect 4387 38165 4399 38168
rect 4341 38159 4399 38165
rect 10042 38156 10048 38168
rect 10100 38156 10106 38208
rect 1104 38106 10856 38128
rect 1104 38054 4213 38106
rect 4265 38054 4277 38106
rect 4329 38054 4341 38106
rect 4393 38054 4405 38106
rect 4457 38054 4469 38106
rect 4521 38054 7477 38106
rect 7529 38054 7541 38106
rect 7593 38054 7605 38106
rect 7657 38054 7669 38106
rect 7721 38054 7733 38106
rect 7785 38054 10856 38106
rect 1104 38032 10856 38054
rect 1394 37952 1400 38004
rect 1452 37992 1458 38004
rect 1489 37995 1547 38001
rect 1489 37992 1501 37995
rect 1452 37964 1501 37992
rect 1452 37952 1458 37964
rect 1489 37961 1501 37964
rect 1535 37961 1547 37995
rect 1489 37955 1547 37961
rect 2501 37995 2559 38001
rect 2501 37961 2513 37995
rect 2547 37992 2559 37995
rect 4062 37992 4068 38004
rect 2547 37964 4068 37992
rect 2547 37961 2559 37964
rect 2501 37955 2559 37961
rect 4062 37952 4068 37964
rect 4120 37952 4126 38004
rect 1854 37924 1860 37936
rect 1504 37896 1860 37924
rect 1504 37800 1532 37896
rect 1854 37884 1860 37896
rect 1912 37884 1918 37936
rect 2314 37924 2320 37936
rect 2148 37896 2320 37924
rect 1673 37859 1731 37865
rect 1673 37825 1685 37859
rect 1719 37856 1731 37859
rect 2148 37856 2176 37896
rect 2314 37884 2320 37896
rect 2372 37884 2378 37936
rect 1719 37828 2176 37856
rect 2225 37859 2283 37865
rect 1719 37825 1731 37828
rect 1673 37819 1731 37825
rect 2225 37825 2237 37859
rect 2271 37825 2283 37859
rect 2498 37856 2504 37868
rect 2459 37828 2504 37856
rect 2225 37819 2283 37825
rect 1486 37748 1492 37800
rect 1544 37748 1550 37800
rect 1854 37748 1860 37800
rect 1912 37788 1918 37800
rect 2240 37788 2268 37819
rect 2498 37816 2504 37828
rect 2556 37816 2562 37868
rect 3053 37859 3111 37865
rect 3053 37825 3065 37859
rect 3099 37856 3111 37859
rect 3694 37856 3700 37868
rect 3099 37828 3700 37856
rect 3099 37825 3111 37828
rect 3053 37819 3111 37825
rect 3694 37816 3700 37828
rect 3752 37816 3758 37868
rect 4154 37856 4160 37868
rect 4115 37828 4160 37856
rect 4154 37816 4160 37828
rect 4212 37816 4218 37868
rect 4341 37859 4399 37865
rect 4341 37825 4353 37859
rect 4387 37856 4399 37859
rect 4614 37856 4620 37868
rect 4387 37828 4620 37856
rect 4387 37825 4399 37828
rect 4341 37819 4399 37825
rect 4614 37816 4620 37828
rect 4672 37816 4678 37868
rect 1912 37760 2268 37788
rect 1912 37748 1918 37760
rect 3234 37652 3240 37664
rect 3195 37624 3240 37652
rect 3234 37612 3240 37624
rect 3292 37612 3298 37664
rect 4341 37655 4399 37661
rect 4341 37621 4353 37655
rect 4387 37652 4399 37655
rect 9858 37652 9864 37664
rect 4387 37624 9864 37652
rect 4387 37621 4399 37624
rect 4341 37615 4399 37621
rect 9858 37612 9864 37624
rect 9916 37612 9922 37664
rect 1104 37562 10856 37584
rect 1104 37510 2582 37562
rect 2634 37510 2646 37562
rect 2698 37510 2710 37562
rect 2762 37510 2774 37562
rect 2826 37510 2838 37562
rect 2890 37510 5845 37562
rect 5897 37510 5909 37562
rect 5961 37510 5973 37562
rect 6025 37510 6037 37562
rect 6089 37510 6101 37562
rect 6153 37510 9109 37562
rect 9161 37510 9173 37562
rect 9225 37510 9237 37562
rect 9289 37510 9301 37562
rect 9353 37510 9365 37562
rect 9417 37510 10856 37562
rect 1104 37488 10856 37510
rect 1486 37272 1492 37324
rect 1544 37272 1550 37324
rect 1397 37247 1455 37253
rect 1397 37213 1409 37247
rect 1443 37244 1455 37247
rect 1504 37244 1532 37272
rect 1443 37216 1532 37244
rect 1443 37213 1455 37216
rect 1397 37207 1455 37213
rect 2038 37204 2044 37256
rect 2096 37244 2102 37256
rect 2133 37247 2191 37253
rect 2133 37244 2145 37247
rect 2096 37216 2145 37244
rect 2096 37204 2102 37216
rect 2133 37213 2145 37216
rect 2179 37213 2191 37247
rect 2958 37244 2964 37256
rect 2919 37216 2964 37244
rect 2133 37207 2191 37213
rect 2958 37204 2964 37216
rect 3016 37204 3022 37256
rect 3053 37247 3111 37253
rect 3053 37213 3065 37247
rect 3099 37244 3111 37247
rect 3786 37244 3792 37256
rect 3099 37216 3792 37244
rect 3099 37213 3111 37216
rect 3053 37207 3111 37213
rect 3786 37204 3792 37216
rect 3844 37204 3850 37256
rect 9858 37244 9864 37256
rect 9819 37216 9864 37244
rect 9858 37204 9864 37216
rect 9916 37204 9922 37256
rect 2406 37136 2412 37188
rect 2464 37176 2470 37188
rect 4154 37176 4160 37188
rect 2464 37148 4160 37176
rect 2464 37136 2470 37148
rect 4154 37136 4160 37148
rect 4212 37136 4218 37188
rect 1578 37108 1584 37120
rect 1539 37080 1584 37108
rect 1578 37068 1584 37080
rect 1636 37068 1642 37120
rect 2314 37108 2320 37120
rect 2275 37080 2320 37108
rect 2314 37068 2320 37080
rect 2372 37068 2378 37120
rect 2958 37068 2964 37120
rect 3016 37108 3022 37120
rect 3142 37108 3148 37120
rect 3016 37080 3148 37108
rect 3016 37068 3022 37080
rect 3142 37068 3148 37080
rect 3200 37068 3206 37120
rect 10042 37108 10048 37120
rect 10003 37080 10048 37108
rect 10042 37068 10048 37080
rect 10100 37068 10106 37120
rect 1104 37018 10856 37040
rect 1104 36966 4213 37018
rect 4265 36966 4277 37018
rect 4329 36966 4341 37018
rect 4393 36966 4405 37018
rect 4457 36966 4469 37018
rect 4521 36966 7477 37018
rect 7529 36966 7541 37018
rect 7593 36966 7605 37018
rect 7657 36966 7669 37018
rect 7721 36966 7733 37018
rect 7785 36966 10856 37018
rect 1104 36944 10856 36966
rect 2225 36907 2283 36913
rect 2225 36873 2237 36907
rect 2271 36904 2283 36907
rect 2406 36904 2412 36916
rect 2271 36876 2412 36904
rect 2271 36873 2283 36876
rect 2225 36867 2283 36873
rect 2406 36864 2412 36876
rect 2464 36864 2470 36916
rect 2869 36907 2927 36913
rect 2869 36873 2881 36907
rect 2915 36904 2927 36907
rect 4798 36904 4804 36916
rect 2915 36876 4804 36904
rect 2915 36873 2927 36876
rect 2869 36867 2927 36873
rect 4798 36864 4804 36876
rect 4856 36864 4862 36916
rect 937 36839 995 36845
rect 937 36805 949 36839
rect 983 36836 995 36839
rect 983 36808 2452 36836
rect 983 36805 995 36808
rect 937 36799 995 36805
rect 2424 36780 2452 36808
rect 1673 36771 1731 36777
rect 1673 36737 1685 36771
rect 1719 36768 1731 36771
rect 1762 36768 1768 36780
rect 1719 36740 1768 36768
rect 1719 36737 1731 36740
rect 1673 36731 1731 36737
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 2038 36728 2044 36780
rect 2096 36768 2102 36780
rect 2317 36771 2375 36777
rect 2317 36768 2329 36771
rect 2096 36740 2329 36768
rect 2096 36728 2102 36740
rect 2317 36737 2329 36740
rect 2363 36737 2375 36771
rect 2317 36731 2375 36737
rect 2406 36728 2412 36780
rect 2464 36728 2470 36780
rect 2777 36771 2835 36777
rect 2777 36737 2789 36771
rect 2823 36768 2835 36771
rect 3510 36768 3516 36780
rect 2823 36740 3516 36768
rect 2823 36737 2835 36740
rect 2777 36731 2835 36737
rect 3510 36728 3516 36740
rect 3568 36728 3574 36780
rect 4157 36771 4215 36777
rect 4157 36737 4169 36771
rect 4203 36737 4215 36771
rect 4157 36731 4215 36737
rect 4341 36771 4399 36777
rect 4341 36737 4353 36771
rect 4387 36768 4399 36771
rect 4614 36768 4620 36780
rect 4387 36740 4620 36768
rect 4387 36737 4399 36740
rect 4341 36731 4399 36737
rect 2222 36660 2228 36712
rect 2280 36700 2286 36712
rect 4172 36700 4200 36731
rect 4614 36728 4620 36740
rect 4672 36728 4678 36780
rect 2280 36672 4200 36700
rect 2280 36660 2286 36672
rect 1486 36564 1492 36576
rect 1447 36536 1492 36564
rect 1486 36524 1492 36536
rect 1544 36524 1550 36576
rect 1670 36524 1676 36576
rect 1728 36564 1734 36576
rect 1854 36564 1860 36576
rect 1728 36536 1860 36564
rect 1728 36524 1734 36536
rect 1854 36524 1860 36536
rect 1912 36524 1918 36576
rect 4341 36567 4399 36573
rect 4341 36533 4353 36567
rect 4387 36564 4399 36567
rect 9858 36564 9864 36576
rect 4387 36536 9864 36564
rect 4387 36533 4399 36536
rect 4341 36527 4399 36533
rect 9858 36524 9864 36536
rect 9916 36524 9922 36576
rect 1104 36474 10856 36496
rect 1104 36422 2582 36474
rect 2634 36422 2646 36474
rect 2698 36422 2710 36474
rect 2762 36422 2774 36474
rect 2826 36422 2838 36474
rect 2890 36422 5845 36474
rect 5897 36422 5909 36474
rect 5961 36422 5973 36474
rect 6025 36422 6037 36474
rect 6089 36422 6101 36474
rect 6153 36422 9109 36474
rect 9161 36422 9173 36474
rect 9225 36422 9237 36474
rect 9289 36422 9301 36474
rect 9353 36422 9365 36474
rect 9417 36422 10856 36474
rect 1104 36400 10856 36422
rect 1394 36320 1400 36372
rect 1452 36360 1458 36372
rect 1670 36360 1676 36372
rect 1452 36332 1676 36360
rect 1452 36320 1458 36332
rect 1670 36320 1676 36332
rect 1728 36320 1734 36372
rect 2222 36360 2228 36372
rect 2183 36332 2228 36360
rect 2222 36320 2228 36332
rect 2280 36320 2286 36372
rect 1397 36159 1455 36165
rect 1397 36125 1409 36159
rect 1443 36156 1455 36159
rect 1946 36156 1952 36168
rect 1443 36128 1952 36156
rect 1443 36125 1455 36128
rect 1397 36119 1455 36125
rect 1946 36116 1952 36128
rect 2004 36116 2010 36168
rect 2222 36116 2228 36168
rect 2280 36156 2286 36168
rect 2317 36159 2375 36165
rect 2317 36156 2329 36159
rect 2280 36128 2329 36156
rect 2280 36116 2286 36128
rect 2317 36125 2329 36128
rect 2363 36125 2375 36159
rect 2317 36119 2375 36125
rect 4157 36159 4215 36165
rect 4157 36125 4169 36159
rect 4203 36125 4215 36159
rect 4157 36119 4215 36125
rect 4341 36159 4399 36165
rect 4341 36125 4353 36159
rect 4387 36156 4399 36159
rect 4614 36156 4620 36168
rect 4387 36128 4620 36156
rect 4387 36125 4399 36128
rect 4341 36119 4399 36125
rect 845 36091 903 36097
rect 845 36057 857 36091
rect 891 36088 903 36091
rect 891 36060 1716 36088
rect 891 36057 903 36060
rect 845 36051 903 36057
rect 1578 36020 1584 36032
rect 1539 35992 1584 36020
rect 1578 35980 1584 35992
rect 1636 35980 1642 36032
rect 1688 36020 1716 36060
rect 1762 36048 1768 36100
rect 1820 36088 1826 36100
rect 4172 36088 4200 36119
rect 4614 36116 4620 36128
rect 4672 36116 4678 36168
rect 9858 36156 9864 36168
rect 9819 36128 9864 36156
rect 9858 36116 9864 36128
rect 9916 36116 9922 36168
rect 1820 36060 4200 36088
rect 1820 36048 1826 36060
rect 1946 36020 1952 36032
rect 1688 35992 1952 36020
rect 1946 35980 1952 35992
rect 2004 35980 2010 36032
rect 4249 36023 4307 36029
rect 4249 35989 4261 36023
rect 4295 36020 4307 36023
rect 9858 36020 9864 36032
rect 4295 35992 9864 36020
rect 4295 35989 4307 35992
rect 4249 35983 4307 35989
rect 9858 35980 9864 35992
rect 9916 35980 9922 36032
rect 10042 36020 10048 36032
rect 10003 35992 10048 36020
rect 10042 35980 10048 35992
rect 10100 35980 10106 36032
rect 1104 35930 10856 35952
rect 1104 35878 4213 35930
rect 4265 35878 4277 35930
rect 4329 35878 4341 35930
rect 4393 35878 4405 35930
rect 4457 35878 4469 35930
rect 4521 35878 7477 35930
rect 7529 35878 7541 35930
rect 7593 35878 7605 35930
rect 7657 35878 7669 35930
rect 7721 35878 7733 35930
rect 7785 35878 10856 35930
rect 1104 35856 10856 35878
rect 2406 35816 2412 35828
rect 2056 35788 2412 35816
rect 1670 35680 1676 35692
rect 1631 35652 1676 35680
rect 1670 35640 1676 35652
rect 1728 35640 1734 35692
rect 2056 35624 2084 35788
rect 2406 35776 2412 35788
rect 2464 35776 2470 35828
rect 2498 35776 2504 35828
rect 2556 35816 2562 35828
rect 2961 35819 3019 35825
rect 2961 35816 2973 35819
rect 2556 35788 2973 35816
rect 2556 35776 2562 35788
rect 2961 35785 2973 35788
rect 3007 35785 3019 35819
rect 2961 35779 3019 35785
rect 3326 35776 3332 35828
rect 3384 35816 3390 35828
rect 3602 35816 3608 35828
rect 3384 35788 3608 35816
rect 3384 35776 3390 35788
rect 3602 35776 3608 35788
rect 3660 35776 3666 35828
rect 2133 35683 2191 35689
rect 2133 35649 2145 35683
rect 2179 35680 2191 35683
rect 2590 35680 2596 35692
rect 2179 35652 2596 35680
rect 2179 35649 2191 35652
rect 2133 35643 2191 35649
rect 2590 35640 2596 35652
rect 2648 35640 2654 35692
rect 3145 35683 3203 35689
rect 3145 35649 3157 35683
rect 3191 35680 3203 35683
rect 3326 35680 3332 35692
rect 3191 35652 3332 35680
rect 3191 35649 3203 35652
rect 3145 35643 3203 35649
rect 3326 35640 3332 35652
rect 3384 35640 3390 35692
rect 2038 35572 2044 35624
rect 2096 35572 2102 35624
rect 2314 35544 2320 35556
rect 2275 35516 2320 35544
rect 2314 35504 2320 35516
rect 2372 35504 2378 35556
rect 1486 35476 1492 35488
rect 1447 35448 1492 35476
rect 1486 35436 1492 35448
rect 1544 35436 1550 35488
rect 1104 35386 10856 35408
rect 1104 35334 2582 35386
rect 2634 35334 2646 35386
rect 2698 35334 2710 35386
rect 2762 35334 2774 35386
rect 2826 35334 2838 35386
rect 2890 35334 5845 35386
rect 5897 35334 5909 35386
rect 5961 35334 5973 35386
rect 6025 35334 6037 35386
rect 6089 35334 6101 35386
rect 6153 35334 9109 35386
rect 9161 35334 9173 35386
rect 9225 35334 9237 35386
rect 9289 35334 9301 35386
rect 9353 35334 9365 35386
rect 9417 35334 10856 35386
rect 1104 35312 10856 35334
rect 4525 35139 4583 35145
rect 4525 35105 4537 35139
rect 4571 35136 4583 35139
rect 4614 35136 4620 35148
rect 4571 35108 4620 35136
rect 4571 35105 4583 35108
rect 4525 35099 4583 35105
rect 4614 35096 4620 35108
rect 4672 35096 4678 35148
rect 1397 35071 1455 35077
rect 1397 35037 1409 35071
rect 1443 35068 1455 35071
rect 1946 35068 1952 35080
rect 1443 35040 1952 35068
rect 1443 35037 1455 35040
rect 1397 35031 1455 35037
rect 1946 35028 1952 35040
rect 2004 35028 2010 35080
rect 4249 35071 4307 35077
rect 4249 35037 4261 35071
rect 4295 35068 4307 35071
rect 4798 35068 4804 35080
rect 4295 35040 4804 35068
rect 4295 35037 4307 35040
rect 4249 35031 4307 35037
rect 4798 35028 4804 35040
rect 4856 35028 4862 35080
rect 9858 35068 9864 35080
rect 9819 35040 9864 35068
rect 9858 35028 9864 35040
rect 9916 35028 9922 35080
rect 1578 34932 1584 34944
rect 1539 34904 1584 34932
rect 1578 34892 1584 34904
rect 1636 34892 1642 34944
rect 1670 34892 1676 34944
rect 1728 34932 1734 34944
rect 3694 34932 3700 34944
rect 1728 34904 3700 34932
rect 1728 34892 1734 34904
rect 3694 34892 3700 34904
rect 3752 34892 3758 34944
rect 10042 34932 10048 34944
rect 10003 34904 10048 34932
rect 10042 34892 10048 34904
rect 10100 34892 10106 34944
rect 1104 34842 10856 34864
rect 1104 34790 4213 34842
rect 4265 34790 4277 34842
rect 4329 34790 4341 34842
rect 4393 34790 4405 34842
rect 4457 34790 4469 34842
rect 4521 34790 7477 34842
rect 7529 34790 7541 34842
rect 7593 34790 7605 34842
rect 7657 34790 7669 34842
rect 7721 34790 7733 34842
rect 7785 34790 10856 34842
rect 1104 34768 10856 34790
rect 2317 34731 2375 34737
rect 2317 34697 2329 34731
rect 2363 34728 2375 34731
rect 5074 34728 5080 34740
rect 2363 34700 5080 34728
rect 2363 34697 2375 34700
rect 2317 34691 2375 34697
rect 5074 34688 5080 34700
rect 5132 34688 5138 34740
rect 3237 34663 3295 34669
rect 3237 34629 3249 34663
rect 3283 34660 3295 34663
rect 5442 34660 5448 34672
rect 3283 34632 5448 34660
rect 3283 34629 3295 34632
rect 3237 34623 3295 34629
rect 5442 34620 5448 34632
rect 5500 34620 5506 34672
rect 1397 34595 1455 34601
rect 1397 34561 1409 34595
rect 1443 34592 1455 34595
rect 1854 34592 1860 34604
rect 1443 34564 1860 34592
rect 1443 34561 1455 34564
rect 1397 34555 1455 34561
rect 1854 34552 1860 34564
rect 1912 34552 1918 34604
rect 2501 34595 2559 34601
rect 2501 34561 2513 34595
rect 2547 34561 2559 34595
rect 3050 34592 3056 34604
rect 3011 34564 3056 34592
rect 2501 34555 2559 34561
rect 2516 34524 2544 34555
rect 3050 34552 3056 34564
rect 3108 34552 3114 34604
rect 3234 34524 3240 34536
rect 2516 34496 3240 34524
rect 3234 34484 3240 34496
rect 3292 34484 3298 34536
rect 1486 34348 1492 34400
rect 1544 34388 1550 34400
rect 1581 34391 1639 34397
rect 1581 34388 1593 34391
rect 1544 34360 1593 34388
rect 1544 34348 1550 34360
rect 1581 34357 1593 34360
rect 1627 34357 1639 34391
rect 1581 34351 1639 34357
rect 1104 34298 10856 34320
rect 1104 34246 2582 34298
rect 2634 34246 2646 34298
rect 2698 34246 2710 34298
rect 2762 34246 2774 34298
rect 2826 34246 2838 34298
rect 2890 34246 5845 34298
rect 5897 34246 5909 34298
rect 5961 34246 5973 34298
rect 6025 34246 6037 34298
rect 6089 34246 6101 34298
rect 6153 34246 9109 34298
rect 9161 34246 9173 34298
rect 9225 34246 9237 34298
rect 9289 34246 9301 34298
rect 9353 34246 9365 34298
rect 9417 34246 10856 34298
rect 1104 34224 10856 34246
rect 3050 34184 3056 34196
rect 3011 34156 3056 34184
rect 3050 34144 3056 34156
rect 3108 34144 3114 34196
rect 1397 33983 1455 33989
rect 1397 33949 1409 33983
rect 1443 33980 1455 33983
rect 2038 33980 2044 33992
rect 1443 33952 2044 33980
rect 1443 33949 1455 33952
rect 1397 33943 1455 33949
rect 2038 33940 2044 33952
rect 2096 33940 2102 33992
rect 2314 33980 2320 33992
rect 2275 33952 2320 33980
rect 2314 33940 2320 33952
rect 2372 33940 2378 33992
rect 2406 33940 2412 33992
rect 2464 33980 2470 33992
rect 2501 33983 2559 33989
rect 2501 33980 2513 33983
rect 2464 33952 2513 33980
rect 2464 33940 2470 33952
rect 2501 33949 2513 33952
rect 2547 33949 2559 33983
rect 2501 33943 2559 33949
rect 3050 33940 3056 33992
rect 3108 33980 3114 33992
rect 3237 33983 3295 33989
rect 3237 33980 3249 33983
rect 3108 33952 3249 33980
rect 3108 33940 3114 33952
rect 3237 33949 3249 33952
rect 3283 33949 3295 33983
rect 9858 33980 9864 33992
rect 9819 33952 9864 33980
rect 3237 33943 3295 33949
rect 9858 33940 9864 33952
rect 9916 33940 9922 33992
rect 7282 33912 7288 33924
rect 2516 33884 7288 33912
rect 1578 33844 1584 33856
rect 1539 33816 1584 33844
rect 1578 33804 1584 33816
rect 1636 33804 1642 33856
rect 2516 33853 2544 33884
rect 7282 33872 7288 33884
rect 7340 33872 7346 33924
rect 2501 33847 2559 33853
rect 2501 33813 2513 33847
rect 2547 33813 2559 33847
rect 2501 33807 2559 33813
rect 2866 33804 2872 33856
rect 2924 33844 2930 33856
rect 5626 33844 5632 33856
rect 2924 33816 5632 33844
rect 2924 33804 2930 33816
rect 5626 33804 5632 33816
rect 5684 33804 5690 33856
rect 10042 33844 10048 33856
rect 10003 33816 10048 33844
rect 10042 33804 10048 33816
rect 10100 33804 10106 33856
rect 1104 33754 10856 33776
rect 1104 33702 4213 33754
rect 4265 33702 4277 33754
rect 4329 33702 4341 33754
rect 4393 33702 4405 33754
rect 4457 33702 4469 33754
rect 4521 33702 7477 33754
rect 7529 33702 7541 33754
rect 7593 33702 7605 33754
rect 7657 33702 7669 33754
rect 7721 33702 7733 33754
rect 7785 33702 10856 33754
rect 1104 33680 10856 33702
rect 2501 33643 2559 33649
rect 2501 33609 2513 33643
rect 2547 33640 2559 33643
rect 2866 33640 2872 33652
rect 2547 33612 2872 33640
rect 2547 33609 2559 33612
rect 2501 33603 2559 33609
rect 2866 33600 2872 33612
rect 2924 33600 2930 33652
rect 3142 33640 3148 33652
rect 3103 33612 3148 33640
rect 3142 33600 3148 33612
rect 3200 33600 3206 33652
rect 2406 33532 2412 33584
rect 2464 33572 2470 33584
rect 2464 33544 4384 33572
rect 2464 33532 2470 33544
rect 1765 33507 1823 33513
rect 1765 33473 1777 33507
rect 1811 33504 1823 33507
rect 2038 33504 2044 33516
rect 1811 33476 2044 33504
rect 1811 33473 1823 33476
rect 1765 33467 1823 33473
rect 2038 33464 2044 33476
rect 2096 33464 2102 33516
rect 2314 33504 2320 33516
rect 2275 33476 2320 33504
rect 2314 33464 2320 33476
rect 2372 33464 2378 33516
rect 2501 33507 2559 33513
rect 2501 33473 2513 33507
rect 2547 33473 2559 33507
rect 3142 33504 3148 33516
rect 3103 33476 3148 33504
rect 2501 33467 2559 33473
rect 1854 33396 1860 33448
rect 1912 33436 1918 33448
rect 2516 33436 2544 33467
rect 3142 33464 3148 33476
rect 3200 33464 3206 33516
rect 3418 33504 3424 33516
rect 3379 33476 3424 33504
rect 3418 33464 3424 33476
rect 3476 33504 3482 33516
rect 4246 33504 4252 33516
rect 3476 33476 4252 33504
rect 3476 33464 3482 33476
rect 4246 33464 4252 33476
rect 4304 33464 4310 33516
rect 4356 33513 4384 33544
rect 4341 33507 4399 33513
rect 4341 33473 4353 33507
rect 4387 33473 4399 33507
rect 4522 33504 4528 33516
rect 4483 33476 4528 33504
rect 4341 33467 4399 33473
rect 4522 33464 4528 33476
rect 4580 33464 4586 33516
rect 1912 33408 2544 33436
rect 1912 33396 1918 33408
rect 4890 33368 4896 33380
rect 3252 33340 4896 33368
rect 1765 33303 1823 33309
rect 1765 33269 1777 33303
rect 1811 33300 1823 33303
rect 3252 33300 3280 33340
rect 4890 33328 4896 33340
rect 4948 33328 4954 33380
rect 1811 33272 3280 33300
rect 4525 33303 4583 33309
rect 1811 33269 1823 33272
rect 1765 33263 1823 33269
rect 4525 33269 4537 33303
rect 4571 33300 4583 33303
rect 9858 33300 9864 33312
rect 4571 33272 9864 33300
rect 4571 33269 4583 33272
rect 4525 33263 4583 33269
rect 9858 33260 9864 33272
rect 9916 33260 9922 33312
rect 1104 33210 10856 33232
rect 1104 33158 2582 33210
rect 2634 33158 2646 33210
rect 2698 33158 2710 33210
rect 2762 33158 2774 33210
rect 2826 33158 2838 33210
rect 2890 33158 5845 33210
rect 5897 33158 5909 33210
rect 5961 33158 5973 33210
rect 6025 33158 6037 33210
rect 6089 33158 6101 33210
rect 6153 33158 9109 33210
rect 9161 33158 9173 33210
rect 9225 33158 9237 33210
rect 9289 33158 9301 33210
rect 9353 33158 9365 33210
rect 9417 33158 10856 33210
rect 1104 33136 10856 33158
rect 3053 33099 3111 33105
rect 3053 33065 3065 33099
rect 3099 33096 3111 33099
rect 3234 33096 3240 33108
rect 3099 33068 3240 33096
rect 3099 33065 3111 33068
rect 3053 33059 3111 33065
rect 3234 33056 3240 33068
rect 3292 33056 3298 33108
rect 1578 33028 1584 33040
rect 1539 33000 1584 33028
rect 1578 32988 1584 33000
rect 1636 32988 1642 33040
rect 2317 33031 2375 33037
rect 2317 32997 2329 33031
rect 2363 33028 2375 33031
rect 5350 33028 5356 33040
rect 2363 33000 5356 33028
rect 2363 32997 2375 33000
rect 2317 32991 2375 32997
rect 5350 32988 5356 33000
rect 5408 32988 5414 33040
rect 2498 32960 2504 32972
rect 1412 32932 2504 32960
rect 1412 32901 1440 32932
rect 2498 32920 2504 32932
rect 2556 32920 2562 32972
rect 1397 32895 1455 32901
rect 1397 32861 1409 32895
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 2314 32852 2320 32904
rect 2372 32892 2378 32904
rect 2409 32895 2467 32901
rect 2409 32892 2421 32895
rect 2372 32864 2421 32892
rect 2372 32852 2378 32864
rect 2409 32861 2421 32864
rect 2455 32861 2467 32895
rect 2409 32855 2467 32861
rect 2593 32895 2651 32901
rect 2593 32861 2605 32895
rect 2639 32892 2651 32895
rect 3234 32892 3240 32904
rect 2639 32864 3004 32892
rect 3195 32864 3240 32892
rect 2639 32861 2651 32864
rect 2593 32855 2651 32861
rect 2424 32824 2452 32855
rect 2774 32824 2780 32836
rect 2424 32796 2780 32824
rect 2774 32784 2780 32796
rect 2832 32784 2838 32836
rect 2976 32824 3004 32864
rect 3234 32852 3240 32864
rect 3292 32852 3298 32904
rect 4246 32852 4252 32904
rect 4304 32892 4310 32904
rect 4341 32895 4399 32901
rect 4341 32892 4353 32895
rect 4304 32864 4353 32892
rect 4304 32852 4310 32864
rect 4341 32861 4353 32864
rect 4387 32861 4399 32895
rect 4522 32892 4528 32904
rect 4483 32864 4528 32892
rect 4341 32855 4399 32861
rect 4522 32852 4528 32864
rect 4580 32852 4586 32904
rect 9861 32895 9919 32901
rect 9861 32892 9873 32895
rect 6886 32864 9873 32892
rect 4890 32824 4896 32836
rect 2976 32796 4896 32824
rect 4890 32784 4896 32796
rect 4948 32784 4954 32836
rect 4433 32759 4491 32765
rect 4433 32725 4445 32759
rect 4479 32756 4491 32759
rect 6886 32756 6914 32864
rect 9861 32861 9873 32864
rect 9907 32861 9919 32895
rect 9861 32855 9919 32861
rect 10042 32756 10048 32768
rect 4479 32728 6914 32756
rect 10003 32728 10048 32756
rect 4479 32725 4491 32728
rect 4433 32719 4491 32725
rect 10042 32716 10048 32728
rect 10100 32716 10106 32768
rect 1104 32666 10856 32688
rect 1104 32614 4213 32666
rect 4265 32614 4277 32666
rect 4329 32614 4341 32666
rect 4393 32614 4405 32666
rect 4457 32614 4469 32666
rect 4521 32614 7477 32666
rect 7529 32614 7541 32666
rect 7593 32614 7605 32666
rect 7657 32614 7669 32666
rect 7721 32614 7733 32666
rect 7785 32614 10856 32666
rect 1104 32592 10856 32614
rect 1581 32555 1639 32561
rect 1581 32521 1593 32555
rect 1627 32552 1639 32555
rect 3510 32552 3516 32564
rect 1627 32524 3516 32552
rect 1627 32521 1639 32524
rect 1581 32515 1639 32521
rect 3510 32512 3516 32524
rect 3568 32512 3574 32564
rect 474 32444 480 32496
rect 532 32484 538 32496
rect 2225 32487 2283 32493
rect 2225 32484 2237 32487
rect 532 32456 2237 32484
rect 532 32444 538 32456
rect 2225 32453 2237 32456
rect 2271 32453 2283 32487
rect 2225 32447 2283 32453
rect 3145 32487 3203 32493
rect 3145 32453 3157 32487
rect 3191 32484 3203 32487
rect 3326 32484 3332 32496
rect 3191 32456 3332 32484
rect 3191 32453 3203 32456
rect 3145 32447 3203 32453
rect 3326 32444 3332 32456
rect 3384 32444 3390 32496
rect 1394 32416 1400 32428
rect 1355 32388 1400 32416
rect 1394 32376 1400 32388
rect 1452 32376 1458 32428
rect 2409 32419 2467 32425
rect 2409 32385 2421 32419
rect 2455 32385 2467 32419
rect 2409 32379 2467 32385
rect 2424 32348 2452 32379
rect 2498 32376 2504 32428
rect 2556 32416 2562 32428
rect 4614 32416 4620 32428
rect 2556 32388 2601 32416
rect 4575 32388 4620 32416
rect 2556 32376 2562 32388
rect 4614 32376 4620 32388
rect 4672 32376 4678 32428
rect 2774 32348 2780 32360
rect 2424 32320 2780 32348
rect 2774 32308 2780 32320
rect 2832 32348 2838 32360
rect 3142 32348 3148 32360
rect 2832 32320 3148 32348
rect 2832 32308 2838 32320
rect 3142 32308 3148 32320
rect 3200 32348 3206 32360
rect 3329 32351 3387 32357
rect 3329 32348 3341 32351
rect 3200 32320 3341 32348
rect 3200 32308 3206 32320
rect 3329 32317 3341 32320
rect 3375 32317 3387 32351
rect 3329 32311 3387 32317
rect 4341 32351 4399 32357
rect 4341 32317 4353 32351
rect 4387 32348 4399 32351
rect 4798 32348 4804 32360
rect 4387 32320 4804 32348
rect 4387 32317 4399 32320
rect 4341 32311 4399 32317
rect 4798 32308 4804 32320
rect 4856 32308 4862 32360
rect 1104 32122 10856 32144
rect 1104 32070 2582 32122
rect 2634 32070 2646 32122
rect 2698 32070 2710 32122
rect 2762 32070 2774 32122
rect 2826 32070 2838 32122
rect 2890 32070 5845 32122
rect 5897 32070 5909 32122
rect 5961 32070 5973 32122
rect 6025 32070 6037 32122
rect 6089 32070 6101 32122
rect 6153 32070 9109 32122
rect 9161 32070 9173 32122
rect 9225 32070 9237 32122
rect 9289 32070 9301 32122
rect 9353 32070 9365 32122
rect 9417 32070 10856 32122
rect 1104 32048 10856 32070
rect 1762 31968 1768 32020
rect 1820 32008 1826 32020
rect 1949 32011 2007 32017
rect 1949 32008 1961 32011
rect 1820 31980 1961 32008
rect 1820 31968 1826 31980
rect 1949 31977 1961 31980
rect 1995 31977 2007 32011
rect 1949 31971 2007 31977
rect 2038 31968 2044 32020
rect 2096 32008 2102 32020
rect 2501 32011 2559 32017
rect 2501 32008 2513 32011
rect 2096 31980 2513 32008
rect 2096 31968 2102 31980
rect 2501 31977 2513 31980
rect 2547 31977 2559 32011
rect 2501 31971 2559 31977
rect 3050 31872 3056 31884
rect 2056 31844 3056 31872
rect 2056 31813 2084 31844
rect 3050 31832 3056 31844
rect 3108 31832 3114 31884
rect 4525 31875 4583 31881
rect 4525 31841 4537 31875
rect 4571 31872 4583 31875
rect 4571 31844 6914 31872
rect 4571 31841 4583 31844
rect 4525 31835 4583 31841
rect 2041 31807 2099 31813
rect 2041 31773 2053 31807
rect 2087 31773 2099 31807
rect 2041 31767 2099 31773
rect 2685 31807 2743 31813
rect 2685 31773 2697 31807
rect 2731 31804 2743 31807
rect 2774 31804 2780 31816
rect 2731 31776 2780 31804
rect 2731 31773 2743 31776
rect 2685 31767 2743 31773
rect 2774 31764 2780 31776
rect 2832 31764 2838 31816
rect 4433 31807 4491 31813
rect 4433 31773 4445 31807
rect 4479 31773 4491 31807
rect 4614 31804 4620 31816
rect 4575 31776 4620 31804
rect 4433 31767 4491 31773
rect 1854 31696 1860 31748
rect 1912 31736 1918 31748
rect 4448 31736 4476 31767
rect 4614 31764 4620 31776
rect 4672 31764 4678 31816
rect 6886 31804 6914 31844
rect 9861 31807 9919 31813
rect 9861 31804 9873 31807
rect 6886 31776 9873 31804
rect 9861 31773 9873 31776
rect 9907 31773 9919 31807
rect 9861 31767 9919 31773
rect 1912 31708 4476 31736
rect 1912 31696 1918 31708
rect 10042 31668 10048 31680
rect 10003 31640 10048 31668
rect 10042 31628 10048 31640
rect 10100 31628 10106 31680
rect 1104 31578 10856 31600
rect 1104 31526 4213 31578
rect 4265 31526 4277 31578
rect 4329 31526 4341 31578
rect 4393 31526 4405 31578
rect 4457 31526 4469 31578
rect 4521 31526 7477 31578
rect 7529 31526 7541 31578
rect 7593 31526 7605 31578
rect 7657 31526 7669 31578
rect 7721 31526 7733 31578
rect 7785 31526 10856 31578
rect 1104 31504 10856 31526
rect 2406 31464 2412 31476
rect 2367 31436 2412 31464
rect 2406 31424 2412 31436
rect 2464 31424 2470 31476
rect 1765 31399 1823 31405
rect 1765 31365 1777 31399
rect 1811 31396 1823 31399
rect 3418 31396 3424 31408
rect 1811 31368 3424 31396
rect 1811 31365 1823 31368
rect 1765 31359 1823 31365
rect 3418 31356 3424 31368
rect 3476 31356 3482 31408
rect 1857 31331 1915 31337
rect 1857 31297 1869 31331
rect 1903 31297 1915 31331
rect 2314 31328 2320 31340
rect 2275 31300 2320 31328
rect 1857 31291 1915 31297
rect 1872 31260 1900 31291
rect 2314 31288 2320 31300
rect 2372 31288 2378 31340
rect 2498 31288 2504 31340
rect 2556 31328 2562 31340
rect 4433 31331 4491 31337
rect 4433 31328 4445 31331
rect 2556 31300 4445 31328
rect 2556 31288 2562 31300
rect 4433 31297 4445 31300
rect 4479 31297 4491 31331
rect 4614 31328 4620 31340
rect 4575 31300 4620 31328
rect 4433 31291 4491 31297
rect 4614 31288 4620 31300
rect 4672 31288 4678 31340
rect 3418 31260 3424 31272
rect 1872 31232 3424 31260
rect 3418 31220 3424 31232
rect 3476 31220 3482 31272
rect 4617 31127 4675 31133
rect 4617 31093 4629 31127
rect 4663 31124 4675 31127
rect 9858 31124 9864 31136
rect 4663 31096 9864 31124
rect 4663 31093 4675 31096
rect 4617 31087 4675 31093
rect 9858 31084 9864 31096
rect 9916 31084 9922 31136
rect 1104 31034 10856 31056
rect 1104 30982 2582 31034
rect 2634 30982 2646 31034
rect 2698 30982 2710 31034
rect 2762 30982 2774 31034
rect 2826 30982 2838 31034
rect 2890 30982 5845 31034
rect 5897 30982 5909 31034
rect 5961 30982 5973 31034
rect 6025 30982 6037 31034
rect 6089 30982 6101 31034
rect 6153 30982 9109 31034
rect 9161 30982 9173 31034
rect 9225 30982 9237 31034
rect 9289 30982 9301 31034
rect 9353 30982 9365 31034
rect 9417 30982 10856 31034
rect 1104 30960 10856 30982
rect 1765 30923 1823 30929
rect 1765 30889 1777 30923
rect 1811 30920 1823 30923
rect 1854 30920 1860 30932
rect 1811 30892 1860 30920
rect 1811 30889 1823 30892
rect 1765 30883 1823 30889
rect 1854 30880 1860 30892
rect 1912 30880 1918 30932
rect 2222 30880 2228 30932
rect 2280 30920 2286 30932
rect 2317 30923 2375 30929
rect 2317 30920 2329 30923
rect 2280 30892 2329 30920
rect 2280 30880 2286 30892
rect 2317 30889 2329 30892
rect 2363 30889 2375 30923
rect 3786 30920 3792 30932
rect 3747 30892 3792 30920
rect 2317 30883 2375 30889
rect 3786 30880 3792 30892
rect 3844 30880 3850 30932
rect 2130 30812 2136 30864
rect 2188 30852 2194 30864
rect 2961 30855 3019 30861
rect 2961 30852 2973 30855
rect 2188 30824 2973 30852
rect 2188 30812 2194 30824
rect 2961 30821 2973 30824
rect 3007 30821 3019 30855
rect 2961 30815 3019 30821
rect 1854 30716 1860 30728
rect 1815 30688 1860 30716
rect 1854 30676 1860 30688
rect 1912 30676 1918 30728
rect 2501 30719 2559 30725
rect 2501 30685 2513 30719
rect 2547 30716 2559 30719
rect 2774 30716 2780 30728
rect 2547 30688 2780 30716
rect 2547 30685 2559 30688
rect 2501 30679 2559 30685
rect 2774 30676 2780 30688
rect 2832 30676 2838 30728
rect 3142 30716 3148 30728
rect 3103 30688 3148 30716
rect 3142 30676 3148 30688
rect 3200 30676 3206 30728
rect 3970 30716 3976 30728
rect 3931 30688 3976 30716
rect 3970 30676 3976 30688
rect 4028 30676 4034 30728
rect 4433 30719 4491 30725
rect 4433 30685 4445 30719
rect 4479 30685 4491 30719
rect 4614 30716 4620 30728
rect 4575 30688 4620 30716
rect 4433 30679 4491 30685
rect 4448 30648 4476 30679
rect 4614 30676 4620 30688
rect 4672 30676 4678 30728
rect 9858 30716 9864 30728
rect 9819 30688 9864 30716
rect 9858 30676 9864 30688
rect 9916 30676 9922 30728
rect 4890 30648 4896 30660
rect 4448 30620 4896 30648
rect 4890 30608 4896 30620
rect 4948 30608 4954 30660
rect 4525 30583 4583 30589
rect 4525 30549 4537 30583
rect 4571 30580 4583 30583
rect 9858 30580 9864 30592
rect 4571 30552 9864 30580
rect 4571 30549 4583 30552
rect 4525 30543 4583 30549
rect 9858 30540 9864 30552
rect 9916 30540 9922 30592
rect 10042 30580 10048 30592
rect 10003 30552 10048 30580
rect 10042 30540 10048 30552
rect 10100 30540 10106 30592
rect 1104 30490 10856 30512
rect 1104 30438 4213 30490
rect 4265 30438 4277 30490
rect 4329 30438 4341 30490
rect 4393 30438 4405 30490
rect 4457 30438 4469 30490
rect 4521 30438 7477 30490
rect 7529 30438 7541 30490
rect 7593 30438 7605 30490
rect 7657 30438 7669 30490
rect 7721 30438 7733 30490
rect 7785 30438 10856 30490
rect 1104 30416 10856 30438
rect 2314 30336 2320 30388
rect 2372 30376 2378 30388
rect 2501 30379 2559 30385
rect 2501 30376 2513 30379
rect 2372 30348 2513 30376
rect 2372 30336 2378 30348
rect 2501 30345 2513 30348
rect 2547 30345 2559 30379
rect 2501 30339 2559 30345
rect 1857 30243 1915 30249
rect 1857 30209 1869 30243
rect 1903 30240 1915 30243
rect 2222 30240 2228 30252
rect 1903 30212 2228 30240
rect 1903 30209 1915 30212
rect 1857 30203 1915 30209
rect 2222 30200 2228 30212
rect 2280 30200 2286 30252
rect 2314 30200 2320 30252
rect 2372 30240 2378 30252
rect 2372 30212 2417 30240
rect 2372 30200 2378 30212
rect 1765 30175 1823 30181
rect 1765 30141 1777 30175
rect 1811 30172 1823 30175
rect 2498 30172 2504 30184
rect 1811 30144 2504 30172
rect 1811 30141 1823 30144
rect 1765 30135 1823 30141
rect 2498 30132 2504 30144
rect 2556 30132 2562 30184
rect 1104 29946 10856 29968
rect 1104 29894 2582 29946
rect 2634 29894 2646 29946
rect 2698 29894 2710 29946
rect 2762 29894 2774 29946
rect 2826 29894 2838 29946
rect 2890 29894 5845 29946
rect 5897 29894 5909 29946
rect 5961 29894 5973 29946
rect 6025 29894 6037 29946
rect 6089 29894 6101 29946
rect 6153 29894 9109 29946
rect 9161 29894 9173 29946
rect 9225 29894 9237 29946
rect 9289 29894 9301 29946
rect 9353 29894 9365 29946
rect 9417 29894 10856 29946
rect 1104 29872 10856 29894
rect 1854 29792 1860 29844
rect 1912 29832 1918 29844
rect 2409 29835 2467 29841
rect 2409 29832 2421 29835
rect 1912 29804 2421 29832
rect 1912 29792 1918 29804
rect 2409 29801 2421 29804
rect 2455 29801 2467 29835
rect 3050 29832 3056 29844
rect 3011 29804 3056 29832
rect 2409 29795 2467 29801
rect 3050 29792 3056 29804
rect 3108 29792 3114 29844
rect 1857 29699 1915 29705
rect 1857 29665 1869 29699
rect 1903 29696 1915 29699
rect 4890 29696 4896 29708
rect 1903 29668 4896 29696
rect 1903 29665 1915 29668
rect 1857 29659 1915 29665
rect 4890 29656 4896 29668
rect 4948 29656 4954 29708
rect 1949 29631 2007 29637
rect 1949 29597 1961 29631
rect 1995 29628 2007 29631
rect 2038 29628 2044 29640
rect 1995 29600 2044 29628
rect 1995 29597 2007 29600
rect 1949 29591 2007 29597
rect 2038 29588 2044 29600
rect 2096 29588 2102 29640
rect 2593 29631 2651 29637
rect 2593 29597 2605 29631
rect 2639 29628 2651 29631
rect 3050 29628 3056 29640
rect 2639 29600 3056 29628
rect 2639 29597 2651 29600
rect 2593 29591 2651 29597
rect 3050 29588 3056 29600
rect 3108 29588 3114 29640
rect 3234 29628 3240 29640
rect 3195 29600 3240 29628
rect 3234 29588 3240 29600
rect 3292 29588 3298 29640
rect 9858 29628 9864 29640
rect 9819 29600 9864 29628
rect 9858 29588 9864 29600
rect 9916 29588 9922 29640
rect 10042 29492 10048 29504
rect 10003 29464 10048 29492
rect 10042 29452 10048 29464
rect 10100 29452 10106 29504
rect 1104 29402 10856 29424
rect 1104 29350 4213 29402
rect 4265 29350 4277 29402
rect 4329 29350 4341 29402
rect 4393 29350 4405 29402
rect 4457 29350 4469 29402
rect 4521 29350 7477 29402
rect 7529 29350 7541 29402
rect 7593 29350 7605 29402
rect 7657 29350 7669 29402
rect 7721 29350 7733 29402
rect 7785 29350 10856 29402
rect 1104 29328 10856 29350
rect 2133 29291 2191 29297
rect 2133 29257 2145 29291
rect 2179 29257 2191 29291
rect 2133 29251 2191 29257
rect 2148 29220 2176 29251
rect 2222 29248 2228 29300
rect 2280 29288 2286 29300
rect 2685 29291 2743 29297
rect 2685 29288 2697 29291
rect 2280 29260 2697 29288
rect 2280 29248 2286 29260
rect 2685 29257 2697 29260
rect 2731 29257 2743 29291
rect 2685 29251 2743 29257
rect 3329 29291 3387 29297
rect 3329 29257 3341 29291
rect 3375 29288 3387 29291
rect 3418 29288 3424 29300
rect 3375 29260 3424 29288
rect 3375 29257 3387 29260
rect 3329 29251 3387 29257
rect 3418 29248 3424 29260
rect 3476 29248 3482 29300
rect 6270 29220 6276 29232
rect 2148 29192 6276 29220
rect 6270 29180 6276 29192
rect 6328 29180 6334 29232
rect 1946 29152 1952 29164
rect 1907 29124 1952 29152
rect 1946 29112 1952 29124
rect 2004 29112 2010 29164
rect 2133 29155 2191 29161
rect 2133 29121 2145 29155
rect 2179 29121 2191 29155
rect 2133 29115 2191 29121
rect 2869 29155 2927 29161
rect 2869 29121 2881 29155
rect 2915 29152 2927 29155
rect 3142 29152 3148 29164
rect 2915 29124 3148 29152
rect 2915 29121 2927 29124
rect 2869 29115 2927 29121
rect 1854 29044 1860 29096
rect 1912 29084 1918 29096
rect 2148 29084 2176 29115
rect 3142 29112 3148 29124
rect 3200 29112 3206 29164
rect 3510 29152 3516 29164
rect 3471 29124 3516 29152
rect 3510 29112 3516 29124
rect 3568 29112 3574 29164
rect 3786 29084 3792 29096
rect 1912 29056 3792 29084
rect 1912 29044 1918 29056
rect 3786 29044 3792 29056
rect 3844 29044 3850 29096
rect 1104 28858 10856 28880
rect 1104 28806 2582 28858
rect 2634 28806 2646 28858
rect 2698 28806 2710 28858
rect 2762 28806 2774 28858
rect 2826 28806 2838 28858
rect 2890 28806 5845 28858
rect 5897 28806 5909 28858
rect 5961 28806 5973 28858
rect 6025 28806 6037 28858
rect 6089 28806 6101 28858
rect 6153 28806 9109 28858
rect 9161 28806 9173 28858
rect 9225 28806 9237 28858
rect 9289 28806 9301 28858
rect 9353 28806 9365 28858
rect 9417 28806 10856 28858
rect 1104 28784 10856 28806
rect 2777 28679 2835 28685
rect 2777 28645 2789 28679
rect 2823 28676 2835 28679
rect 3602 28676 3608 28688
rect 2823 28648 3608 28676
rect 2823 28645 2835 28648
rect 2777 28639 2835 28645
rect 3602 28636 3608 28648
rect 3660 28636 3666 28688
rect 566 28568 572 28620
rect 624 28608 630 28620
rect 1857 28611 1915 28617
rect 1857 28608 1869 28611
rect 624 28580 1869 28608
rect 624 28568 630 28580
rect 1857 28577 1869 28580
rect 1903 28577 1915 28611
rect 1857 28571 1915 28577
rect 1946 28500 1952 28552
rect 2004 28540 2010 28552
rect 2041 28543 2099 28549
rect 2041 28540 2053 28543
rect 2004 28512 2053 28540
rect 2004 28500 2010 28512
rect 2041 28509 2053 28512
rect 2087 28509 2099 28543
rect 2041 28503 2099 28509
rect 2056 28472 2084 28503
rect 2130 28500 2136 28552
rect 2188 28540 2194 28552
rect 2866 28540 2872 28552
rect 2188 28512 2233 28540
rect 2827 28512 2872 28540
rect 2188 28500 2194 28512
rect 2866 28500 2872 28512
rect 2924 28500 2930 28552
rect 3053 28543 3111 28549
rect 3053 28509 3065 28543
rect 3099 28540 3111 28543
rect 3694 28540 3700 28552
rect 3099 28512 3700 28540
rect 3099 28509 3111 28512
rect 3053 28503 3111 28509
rect 3694 28500 3700 28512
rect 3752 28500 3758 28552
rect 3786 28500 3792 28552
rect 3844 28540 3850 28552
rect 3973 28543 4031 28549
rect 3844 28512 3889 28540
rect 3844 28500 3850 28512
rect 3973 28509 3985 28543
rect 4019 28540 4031 28543
rect 4614 28540 4620 28552
rect 4019 28512 4620 28540
rect 4019 28509 4031 28512
rect 3973 28503 4031 28509
rect 4614 28500 4620 28512
rect 4672 28500 4678 28552
rect 9861 28543 9919 28549
rect 9861 28540 9873 28543
rect 6886 28512 9873 28540
rect 2884 28472 2912 28500
rect 2056 28444 2912 28472
rect 3881 28407 3939 28413
rect 3881 28373 3893 28407
rect 3927 28404 3939 28407
rect 6886 28404 6914 28512
rect 9861 28509 9873 28512
rect 9907 28509 9919 28543
rect 9861 28503 9919 28509
rect 10042 28404 10048 28416
rect 3927 28376 6914 28404
rect 10003 28376 10048 28404
rect 3927 28373 3939 28376
rect 3881 28367 3939 28373
rect 10042 28364 10048 28376
rect 10100 28364 10106 28416
rect 1104 28314 10856 28336
rect 1104 28262 4213 28314
rect 4265 28262 4277 28314
rect 4329 28262 4341 28314
rect 4393 28262 4405 28314
rect 4457 28262 4469 28314
rect 4521 28262 7477 28314
rect 7529 28262 7541 28314
rect 7593 28262 7605 28314
rect 7657 28262 7669 28314
rect 7721 28262 7733 28314
rect 7785 28262 10856 28314
rect 1104 28240 10856 28262
rect 2958 28200 2964 28212
rect 2919 28172 2964 28200
rect 2958 28160 2964 28172
rect 3016 28160 3022 28212
rect 2225 28135 2283 28141
rect 2225 28101 2237 28135
rect 2271 28132 2283 28135
rect 6178 28132 6184 28144
rect 2271 28104 6184 28132
rect 2271 28101 2283 28104
rect 2225 28095 2283 28101
rect 6178 28092 6184 28104
rect 6236 28092 6242 28144
rect 1486 28024 1492 28076
rect 1544 28064 1550 28076
rect 1857 28067 1915 28073
rect 1857 28064 1869 28067
rect 1544 28036 1869 28064
rect 1544 28024 1550 28036
rect 1857 28033 1869 28036
rect 1903 28033 1915 28067
rect 1857 28027 1915 28033
rect 2133 28067 2191 28073
rect 2133 28033 2145 28067
rect 2179 28064 2191 28067
rect 2866 28064 2872 28076
rect 2179 28036 2872 28064
rect 2179 28033 2191 28036
rect 2133 28027 2191 28033
rect 2866 28024 2872 28036
rect 2924 28024 2930 28076
rect 3053 28067 3111 28073
rect 3053 28033 3065 28067
rect 3099 28064 3111 28067
rect 3234 28064 3240 28076
rect 3099 28036 3240 28064
rect 3099 28033 3111 28036
rect 3053 28027 3111 28033
rect 3234 28024 3240 28036
rect 3292 28024 3298 28076
rect 3973 28067 4031 28073
rect 3973 28033 3985 28067
rect 4019 28064 4031 28067
rect 4522 28064 4528 28076
rect 4019 28036 4528 28064
rect 4019 28033 4031 28036
rect 3973 28027 4031 28033
rect 4522 28024 4528 28036
rect 4580 28064 4586 28076
rect 4798 28064 4804 28076
rect 4580 28036 4804 28064
rect 4580 28024 4586 28036
rect 4798 28024 4804 28036
rect 4856 28024 4862 28076
rect 4246 27996 4252 28008
rect 4207 27968 4252 27996
rect 4246 27956 4252 27968
rect 4304 27996 4310 28008
rect 4614 27996 4620 28008
rect 4304 27968 4620 27996
rect 4304 27956 4310 27968
rect 4614 27956 4620 27968
rect 4672 27956 4678 28008
rect 1104 27770 10856 27792
rect 1104 27718 2582 27770
rect 2634 27718 2646 27770
rect 2698 27718 2710 27770
rect 2762 27718 2774 27770
rect 2826 27718 2838 27770
rect 2890 27718 5845 27770
rect 5897 27718 5909 27770
rect 5961 27718 5973 27770
rect 6025 27718 6037 27770
rect 6089 27718 6101 27770
rect 6153 27718 9109 27770
rect 9161 27718 9173 27770
rect 9225 27718 9237 27770
rect 9289 27718 9301 27770
rect 9353 27718 9365 27770
rect 9417 27718 10856 27770
rect 1104 27696 10856 27718
rect 2869 27659 2927 27665
rect 2869 27625 2881 27659
rect 2915 27656 2927 27659
rect 2958 27656 2964 27668
rect 2915 27628 2964 27656
rect 2915 27625 2927 27628
rect 2869 27619 2927 27625
rect 2958 27616 2964 27628
rect 3016 27616 3022 27668
rect 1489 27591 1547 27597
rect 1489 27557 1501 27591
rect 1535 27588 1547 27591
rect 1854 27588 1860 27600
rect 1535 27560 1860 27588
rect 1535 27557 1547 27560
rect 1489 27551 1547 27557
rect 1854 27548 1860 27560
rect 1912 27548 1918 27600
rect 2038 27588 2044 27600
rect 1999 27560 2044 27588
rect 2038 27548 2044 27560
rect 2096 27548 2102 27600
rect 1578 27452 1584 27464
rect 1539 27424 1584 27452
rect 1578 27412 1584 27424
rect 1636 27412 1642 27464
rect 2222 27452 2228 27464
rect 2183 27424 2228 27452
rect 2222 27412 2228 27424
rect 2280 27412 2286 27464
rect 2961 27455 3019 27461
rect 2961 27421 2973 27455
rect 3007 27452 3019 27455
rect 3050 27452 3056 27464
rect 3007 27424 3056 27452
rect 3007 27421 3019 27424
rect 2961 27415 3019 27421
rect 3050 27412 3056 27424
rect 3108 27452 3114 27464
rect 3326 27452 3332 27464
rect 3108 27424 3332 27452
rect 3108 27412 3114 27424
rect 3326 27412 3332 27424
rect 3384 27412 3390 27464
rect 3694 27412 3700 27464
rect 3752 27452 3758 27464
rect 3789 27455 3847 27461
rect 3789 27452 3801 27455
rect 3752 27424 3801 27452
rect 3752 27412 3758 27424
rect 3789 27421 3801 27424
rect 3835 27421 3847 27455
rect 3970 27452 3976 27464
rect 3931 27424 3976 27452
rect 3789 27415 3847 27421
rect 3970 27412 3976 27424
rect 4028 27452 4034 27464
rect 4246 27452 4252 27464
rect 4028 27424 4252 27452
rect 4028 27412 4034 27424
rect 4246 27412 4252 27424
rect 4304 27412 4310 27464
rect 9861 27455 9919 27461
rect 9861 27452 9873 27455
rect 6886 27424 9873 27452
rect 3881 27319 3939 27325
rect 3881 27285 3893 27319
rect 3927 27316 3939 27319
rect 6886 27316 6914 27424
rect 9861 27421 9873 27424
rect 9907 27421 9919 27455
rect 9861 27415 9919 27421
rect 10042 27316 10048 27328
rect 3927 27288 6914 27316
rect 10003 27288 10048 27316
rect 3927 27285 3939 27288
rect 3881 27279 3939 27285
rect 10042 27276 10048 27288
rect 10100 27276 10106 27328
rect 1104 27226 10856 27248
rect 1104 27174 4213 27226
rect 4265 27174 4277 27226
rect 4329 27174 4341 27226
rect 4393 27174 4405 27226
rect 4457 27174 4469 27226
rect 4521 27174 7477 27226
rect 7529 27174 7541 27226
rect 7593 27174 7605 27226
rect 7657 27174 7669 27226
rect 7721 27174 7733 27226
rect 7785 27174 10856 27226
rect 1104 27152 10856 27174
rect 1578 27072 1584 27124
rect 1636 27112 1642 27124
rect 2685 27115 2743 27121
rect 2685 27112 2697 27115
rect 1636 27084 2697 27112
rect 1636 27072 1642 27084
rect 2685 27081 2697 27084
rect 2731 27081 2743 27115
rect 2685 27075 2743 27081
rect 2133 27047 2191 27053
rect 2133 27013 2145 27047
rect 2179 27044 2191 27047
rect 3694 27044 3700 27056
rect 2179 27016 3700 27044
rect 2179 27013 2191 27016
rect 2133 27007 2191 27013
rect 3694 27004 3700 27016
rect 3752 27004 3758 27056
rect 1578 26976 1584 26988
rect 1539 26948 1584 26976
rect 1578 26936 1584 26948
rect 1636 26936 1642 26988
rect 2041 26979 2099 26985
rect 2041 26945 2053 26979
rect 2087 26976 2099 26979
rect 2222 26976 2228 26988
rect 2087 26948 2228 26976
rect 2087 26945 2099 26948
rect 2041 26939 2099 26945
rect 2222 26936 2228 26948
rect 2280 26936 2286 26988
rect 2866 26976 2872 26988
rect 2827 26948 2872 26976
rect 2866 26936 2872 26948
rect 2924 26936 2930 26988
rect 3605 26979 3663 26985
rect 3605 26945 3617 26979
rect 3651 26945 3663 26979
rect 3605 26939 3663 26945
rect 3789 26979 3847 26985
rect 3789 26945 3801 26979
rect 3835 26976 3847 26979
rect 3970 26976 3976 26988
rect 3835 26948 3976 26976
rect 3835 26945 3847 26948
rect 3789 26939 3847 26945
rect 1489 26911 1547 26917
rect 1489 26877 1501 26911
rect 1535 26908 1547 26911
rect 2130 26908 2136 26920
rect 1535 26880 2136 26908
rect 1535 26877 1547 26880
rect 1489 26871 1547 26877
rect 2130 26868 2136 26880
rect 2188 26908 2194 26920
rect 3620 26908 3648 26939
rect 3970 26936 3976 26948
rect 4028 26976 4034 26988
rect 4154 26976 4160 26988
rect 4028 26948 4160 26976
rect 4028 26936 4034 26948
rect 4154 26936 4160 26948
rect 4212 26936 4218 26988
rect 2188 26880 3648 26908
rect 2188 26868 2194 26880
rect 3789 26775 3847 26781
rect 3789 26741 3801 26775
rect 3835 26772 3847 26775
rect 9858 26772 9864 26784
rect 3835 26744 9864 26772
rect 3835 26741 3847 26744
rect 3789 26735 3847 26741
rect 9858 26732 9864 26744
rect 9916 26732 9922 26784
rect 1104 26682 10856 26704
rect 1104 26630 2582 26682
rect 2634 26630 2646 26682
rect 2698 26630 2710 26682
rect 2762 26630 2774 26682
rect 2826 26630 2838 26682
rect 2890 26630 5845 26682
rect 5897 26630 5909 26682
rect 5961 26630 5973 26682
rect 6025 26630 6037 26682
rect 6089 26630 6101 26682
rect 6153 26630 9109 26682
rect 9161 26630 9173 26682
rect 9225 26630 9237 26682
rect 9289 26630 9301 26682
rect 9353 26630 9365 26682
rect 9417 26630 10856 26682
rect 1104 26608 10856 26630
rect 2222 26568 2228 26580
rect 2183 26540 2228 26568
rect 2222 26528 2228 26540
rect 2280 26528 2286 26580
rect 3973 26571 4031 26577
rect 3973 26537 3985 26571
rect 4019 26568 4031 26571
rect 4019 26540 4568 26568
rect 4019 26537 4031 26540
rect 3973 26531 4031 26537
rect 1489 26503 1547 26509
rect 1489 26469 1501 26503
rect 1535 26500 1547 26503
rect 3234 26500 3240 26512
rect 1535 26472 3240 26500
rect 1535 26469 1547 26472
rect 1489 26463 1547 26469
rect 3234 26460 3240 26472
rect 3292 26500 3298 26512
rect 3292 26472 4476 26500
rect 3292 26460 3298 26472
rect 658 26392 664 26444
rect 716 26432 722 26444
rect 2869 26435 2927 26441
rect 2869 26432 2881 26435
rect 716 26404 2881 26432
rect 716 26392 722 26404
rect 2869 26401 2881 26404
rect 2915 26401 2927 26435
rect 2869 26395 2927 26401
rect 1581 26367 1639 26373
rect 1581 26333 1593 26367
rect 1627 26364 1639 26367
rect 1854 26364 1860 26376
rect 1627 26336 1860 26364
rect 1627 26333 1639 26336
rect 1581 26327 1639 26333
rect 1854 26324 1860 26336
rect 1912 26324 1918 26376
rect 2038 26364 2044 26376
rect 1999 26336 2044 26364
rect 2038 26324 2044 26336
rect 2096 26324 2102 26376
rect 3786 26364 3792 26376
rect 3747 26336 3792 26364
rect 3786 26324 3792 26336
rect 3844 26324 3850 26376
rect 4448 26373 4476 26472
rect 4540 26432 4568 26540
rect 4617 26503 4675 26509
rect 4617 26469 4629 26503
rect 4663 26500 4675 26503
rect 9950 26500 9956 26512
rect 4663 26472 9956 26500
rect 4663 26469 4675 26472
rect 4617 26463 4675 26469
rect 9950 26460 9956 26472
rect 10008 26460 10014 26512
rect 4540 26404 5396 26432
rect 3973 26367 4031 26373
rect 3973 26333 3985 26367
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4433 26367 4491 26373
rect 4433 26333 4445 26367
rect 4479 26333 4491 26367
rect 4433 26327 4491 26333
rect 4617 26367 4675 26373
rect 4617 26333 4629 26367
rect 4663 26333 4675 26367
rect 4617 26327 4675 26333
rect 3145 26299 3203 26305
rect 3145 26265 3157 26299
rect 3191 26296 3203 26299
rect 3234 26296 3240 26308
rect 3191 26268 3240 26296
rect 3191 26265 3203 26268
rect 3145 26259 3203 26265
rect 3234 26256 3240 26268
rect 3292 26256 3298 26308
rect 3988 26296 4016 26327
rect 4154 26296 4160 26308
rect 3988 26268 4160 26296
rect 4154 26256 4160 26268
rect 4212 26296 4218 26308
rect 4632 26296 4660 26327
rect 4212 26268 4660 26296
rect 5368 26296 5396 26404
rect 9858 26364 9864 26376
rect 9819 26336 9864 26364
rect 9858 26324 9864 26336
rect 9916 26324 9922 26376
rect 9766 26296 9772 26308
rect 5368 26268 9772 26296
rect 4212 26256 4218 26268
rect 9766 26256 9772 26268
rect 9824 26256 9830 26308
rect 1486 26188 1492 26240
rect 1544 26228 1550 26240
rect 3786 26228 3792 26240
rect 1544 26200 3792 26228
rect 1544 26188 1550 26200
rect 3786 26188 3792 26200
rect 3844 26188 3850 26240
rect 10042 26228 10048 26240
rect 10003 26200 10048 26228
rect 10042 26188 10048 26200
rect 10100 26188 10106 26240
rect 1104 26138 10856 26160
rect 1104 26086 4213 26138
rect 4265 26086 4277 26138
rect 4329 26086 4341 26138
rect 4393 26086 4405 26138
rect 4457 26086 4469 26138
rect 4521 26086 7477 26138
rect 7529 26086 7541 26138
rect 7593 26086 7605 26138
rect 7657 26086 7669 26138
rect 7721 26086 7733 26138
rect 7785 26086 10856 26138
rect 1104 26064 10856 26086
rect 1486 26024 1492 26036
rect 1447 25996 1492 26024
rect 1486 25984 1492 25996
rect 1544 25984 1550 26036
rect 1578 25984 1584 26036
rect 1636 26024 1642 26036
rect 2041 26027 2099 26033
rect 2041 26024 2053 26027
rect 1636 25996 2053 26024
rect 1636 25984 1642 25996
rect 2041 25993 2053 25996
rect 2087 25993 2099 26027
rect 2041 25987 2099 25993
rect 1581 25891 1639 25897
rect 1581 25857 1593 25891
rect 1627 25888 1639 25891
rect 2038 25888 2044 25900
rect 1627 25860 2044 25888
rect 1627 25857 1639 25860
rect 1581 25851 1639 25857
rect 2038 25848 2044 25860
rect 2096 25848 2102 25900
rect 2222 25888 2228 25900
rect 2183 25860 2228 25888
rect 2222 25848 2228 25860
rect 2280 25848 2286 25900
rect 1104 25594 10856 25616
rect 1104 25542 2582 25594
rect 2634 25542 2646 25594
rect 2698 25542 2710 25594
rect 2762 25542 2774 25594
rect 2826 25542 2838 25594
rect 2890 25542 5845 25594
rect 5897 25542 5909 25594
rect 5961 25542 5973 25594
rect 6025 25542 6037 25594
rect 6089 25542 6101 25594
rect 6153 25542 9109 25594
rect 9161 25542 9173 25594
rect 9225 25542 9237 25594
rect 9289 25542 9301 25594
rect 9353 25542 9365 25594
rect 9417 25542 10856 25594
rect 1104 25520 10856 25542
rect 2038 25480 2044 25492
rect 1999 25452 2044 25480
rect 2038 25440 2044 25452
rect 2096 25440 2102 25492
rect 1854 25372 1860 25424
rect 1912 25412 1918 25424
rect 2685 25415 2743 25421
rect 2685 25412 2697 25415
rect 1912 25384 2697 25412
rect 1912 25372 1918 25384
rect 2685 25381 2697 25384
rect 2731 25381 2743 25415
rect 2685 25375 2743 25381
rect 4062 25304 4068 25356
rect 4120 25344 4126 25356
rect 6362 25344 6368 25356
rect 4120 25316 6368 25344
rect 4120 25304 4126 25316
rect 6362 25304 6368 25316
rect 6420 25304 6426 25356
rect 1394 25276 1400 25288
rect 1355 25248 1400 25276
rect 1394 25236 1400 25248
rect 1452 25236 1458 25288
rect 2222 25276 2228 25288
rect 2183 25248 2228 25276
rect 2222 25236 2228 25248
rect 2280 25236 2286 25288
rect 2866 25276 2872 25288
rect 2827 25248 2872 25276
rect 2866 25236 2872 25248
rect 2924 25236 2930 25288
rect 9861 25279 9919 25285
rect 9861 25245 9873 25279
rect 9907 25276 9919 25279
rect 9950 25276 9956 25288
rect 9907 25248 9956 25276
rect 9907 25245 9919 25248
rect 9861 25239 9919 25245
rect 9950 25236 9956 25248
rect 10008 25236 10014 25288
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 2038 25140 2044 25152
rect 1627 25112 2044 25140
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 2038 25100 2044 25112
rect 2096 25100 2102 25152
rect 10042 25140 10048 25152
rect 10003 25112 10048 25140
rect 10042 25100 10048 25112
rect 10100 25100 10106 25152
rect 1104 25050 10856 25072
rect 1104 24998 4213 25050
rect 4265 24998 4277 25050
rect 4329 24998 4341 25050
rect 4393 24998 4405 25050
rect 4457 24998 4469 25050
rect 4521 24998 7477 25050
rect 7529 24998 7541 25050
rect 7593 24998 7605 25050
rect 7657 24998 7669 25050
rect 7721 24998 7733 25050
rect 7785 24998 10856 25050
rect 1104 24976 10856 24998
rect 1397 24803 1455 24809
rect 1397 24769 1409 24803
rect 1443 24800 1455 24803
rect 1486 24800 1492 24812
rect 1443 24772 1492 24800
rect 1443 24769 1455 24772
rect 1397 24763 1455 24769
rect 1486 24760 1492 24772
rect 1544 24760 1550 24812
rect 3234 24800 3240 24812
rect 3195 24772 3240 24800
rect 3234 24760 3240 24772
rect 3292 24760 3298 24812
rect 3329 24803 3387 24809
rect 3329 24769 3341 24803
rect 3375 24800 3387 24803
rect 4065 24803 4123 24809
rect 4065 24800 4077 24803
rect 3375 24772 4077 24800
rect 3375 24769 3387 24772
rect 3329 24763 3387 24769
rect 4065 24769 4077 24772
rect 4111 24800 4123 24803
rect 4246 24800 4252 24812
rect 4111 24772 4252 24800
rect 4111 24769 4123 24772
rect 4065 24763 4123 24769
rect 4246 24760 4252 24772
rect 4304 24760 4310 24812
rect 1394 24556 1400 24608
rect 1452 24596 1458 24608
rect 1581 24599 1639 24605
rect 1581 24596 1593 24599
rect 1452 24568 1593 24596
rect 1452 24556 1458 24568
rect 1581 24565 1593 24568
rect 1627 24565 1639 24599
rect 1581 24559 1639 24565
rect 4341 24599 4399 24605
rect 4341 24565 4353 24599
rect 4387 24596 4399 24599
rect 4982 24596 4988 24608
rect 4387 24568 4988 24596
rect 4387 24565 4399 24568
rect 4341 24559 4399 24565
rect 4982 24556 4988 24568
rect 5040 24556 5046 24608
rect 1104 24506 10856 24528
rect 1104 24454 2582 24506
rect 2634 24454 2646 24506
rect 2698 24454 2710 24506
rect 2762 24454 2774 24506
rect 2826 24454 2838 24506
rect 2890 24454 5845 24506
rect 5897 24454 5909 24506
rect 5961 24454 5973 24506
rect 6025 24454 6037 24506
rect 6089 24454 6101 24506
rect 6153 24454 9109 24506
rect 9161 24454 9173 24506
rect 9225 24454 9237 24506
rect 9289 24454 9301 24506
rect 9353 24454 9365 24506
rect 9417 24454 10856 24506
rect 1104 24432 10856 24454
rect 3878 24352 3884 24404
rect 3936 24392 3942 24404
rect 4706 24392 4712 24404
rect 3936 24364 4712 24392
rect 3936 24352 3942 24364
rect 4706 24352 4712 24364
rect 4764 24352 4770 24404
rect 2685 24327 2743 24333
rect 2685 24293 2697 24327
rect 2731 24293 2743 24327
rect 2685 24287 2743 24293
rect 4433 24327 4491 24333
rect 4433 24293 4445 24327
rect 4479 24324 4491 24327
rect 4614 24324 4620 24336
rect 4479 24296 4620 24324
rect 4479 24293 4491 24296
rect 4433 24287 4491 24293
rect 2700 24256 2728 24287
rect 4614 24284 4620 24296
rect 4672 24284 4678 24336
rect 1596 24228 2728 24256
rect 1596 24197 1624 24228
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24157 1639 24191
rect 2038 24188 2044 24200
rect 1999 24160 2044 24188
rect 1581 24151 1639 24157
rect 2038 24148 2044 24160
rect 2096 24148 2102 24200
rect 2866 24188 2872 24200
rect 2827 24160 2872 24188
rect 2866 24148 2872 24160
rect 2924 24148 2930 24200
rect 4246 24188 4252 24200
rect 4207 24160 4252 24188
rect 4246 24148 4252 24160
rect 4304 24148 4310 24200
rect 9766 24148 9772 24200
rect 9824 24188 9830 24200
rect 9861 24191 9919 24197
rect 9861 24188 9873 24191
rect 9824 24160 9873 24188
rect 9824 24148 9830 24160
rect 9861 24157 9873 24160
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 1489 24055 1547 24061
rect 1489 24021 1501 24055
rect 1535 24052 1547 24055
rect 2038 24052 2044 24064
rect 1535 24024 2044 24052
rect 1535 24021 1547 24024
rect 1489 24015 1547 24021
rect 2038 24012 2044 24024
rect 2096 24012 2102 24064
rect 2130 24012 2136 24064
rect 2188 24052 2194 24064
rect 10042 24052 10048 24064
rect 2188 24024 2233 24052
rect 10003 24024 10048 24052
rect 2188 24012 2194 24024
rect 10042 24012 10048 24024
rect 10100 24012 10106 24064
rect 1104 23962 10856 23984
rect 1104 23910 4213 23962
rect 4265 23910 4277 23962
rect 4329 23910 4341 23962
rect 4393 23910 4405 23962
rect 4457 23910 4469 23962
rect 4521 23910 7477 23962
rect 7529 23910 7541 23962
rect 7593 23910 7605 23962
rect 7657 23910 7669 23962
rect 7721 23910 7733 23962
rect 7785 23910 10856 23962
rect 1104 23888 10856 23910
rect 3053 23851 3111 23857
rect 3053 23817 3065 23851
rect 3099 23848 3111 23851
rect 4062 23848 4068 23860
rect 3099 23820 4068 23848
rect 3099 23817 3111 23820
rect 3053 23811 3111 23817
rect 4062 23808 4068 23820
rect 4120 23808 4126 23860
rect 2130 23740 2136 23792
rect 2188 23780 2194 23792
rect 4338 23780 4344 23792
rect 2188 23752 4344 23780
rect 2188 23740 2194 23752
rect 2038 23712 2044 23724
rect 1951 23684 2044 23712
rect 2038 23672 2044 23684
rect 2096 23672 2102 23724
rect 2225 23715 2283 23721
rect 2225 23681 2237 23715
rect 2271 23712 2283 23715
rect 2958 23712 2964 23724
rect 2271 23684 2964 23712
rect 2271 23681 2283 23684
rect 2225 23675 2283 23681
rect 2958 23672 2964 23684
rect 3016 23672 3022 23724
rect 3160 23721 3188 23752
rect 4338 23740 4344 23752
rect 4396 23740 4402 23792
rect 3145 23715 3203 23721
rect 3145 23681 3157 23715
rect 3191 23681 3203 23715
rect 3786 23712 3792 23724
rect 3747 23684 3792 23712
rect 3145 23675 3203 23681
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 2056 23644 2084 23672
rect 4062 23644 4068 23656
rect 2056 23616 4068 23644
rect 4062 23604 4068 23616
rect 4120 23604 4126 23656
rect 2225 23579 2283 23585
rect 2225 23545 2237 23579
rect 2271 23576 2283 23579
rect 6546 23576 6552 23588
rect 2271 23548 6552 23576
rect 2271 23545 2283 23548
rect 2225 23539 2283 23545
rect 6546 23536 6552 23548
rect 6604 23536 6610 23588
rect 3602 23508 3608 23520
rect 3563 23480 3608 23508
rect 3602 23468 3608 23480
rect 3660 23468 3666 23520
rect 1104 23418 10856 23440
rect 1104 23366 2582 23418
rect 2634 23366 2646 23418
rect 2698 23366 2710 23418
rect 2762 23366 2774 23418
rect 2826 23366 2838 23418
rect 2890 23366 5845 23418
rect 5897 23366 5909 23418
rect 5961 23366 5973 23418
rect 6025 23366 6037 23418
rect 6089 23366 6101 23418
rect 6153 23366 9109 23418
rect 9161 23366 9173 23418
rect 9225 23366 9237 23418
rect 9289 23366 9301 23418
rect 9353 23366 9365 23418
rect 9417 23366 10856 23418
rect 1104 23344 10856 23366
rect 3050 23304 3056 23316
rect 3011 23276 3056 23304
rect 3050 23264 3056 23276
rect 3108 23264 3114 23316
rect 2038 23168 2044 23180
rect 1999 23140 2044 23168
rect 2038 23128 2044 23140
rect 2096 23128 2102 23180
rect 2958 23168 2964 23180
rect 2240 23140 2964 23168
rect 1394 23100 1400 23112
rect 1355 23072 1400 23100
rect 1394 23060 1400 23072
rect 1452 23060 1458 23112
rect 2240 23109 2268 23140
rect 2958 23128 2964 23140
rect 3016 23128 3022 23180
rect 4614 23168 4620 23180
rect 4264 23140 4620 23168
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23069 2283 23103
rect 2225 23063 2283 23069
rect 2409 23103 2467 23109
rect 2409 23069 2421 23103
rect 2455 23100 2467 23103
rect 3142 23100 3148 23112
rect 2455 23072 3148 23100
rect 2455 23069 2467 23072
rect 2409 23063 2467 23069
rect 1489 23035 1547 23041
rect 1489 23001 1501 23035
rect 1535 23032 1547 23035
rect 2424 23032 2452 23063
rect 3142 23060 3148 23072
rect 3200 23060 3206 23112
rect 4062 23100 4068 23112
rect 4023 23072 4068 23100
rect 4062 23060 4068 23072
rect 4120 23060 4126 23112
rect 4264 23109 4292 23140
rect 4614 23128 4620 23140
rect 4672 23168 4678 23180
rect 4672 23140 4936 23168
rect 4672 23128 4678 23140
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23069 4307 23103
rect 4249 23063 4307 23069
rect 4338 23060 4344 23112
rect 4396 23100 4402 23112
rect 4908 23109 4936 23140
rect 4709 23103 4767 23109
rect 4709 23100 4721 23103
rect 4396 23072 4721 23100
rect 4396 23060 4402 23072
rect 4709 23069 4721 23072
rect 4755 23069 4767 23103
rect 4709 23063 4767 23069
rect 4893 23103 4951 23109
rect 4893 23069 4905 23103
rect 4939 23069 4951 23103
rect 9861 23103 9919 23109
rect 9861 23100 9873 23103
rect 4893 23063 4951 23069
rect 6886 23072 9873 23100
rect 1535 23004 2452 23032
rect 2961 23035 3019 23041
rect 1535 23001 1547 23004
rect 1489 22995 1547 23001
rect 2961 23001 2973 23035
rect 3007 23032 3019 23035
rect 3418 23032 3424 23044
rect 3007 23004 3424 23032
rect 3007 23001 3019 23004
rect 2961 22995 3019 23001
rect 3418 22992 3424 23004
rect 3476 23032 3482 23044
rect 6638 23032 6644 23044
rect 3476 23004 6644 23032
rect 3476 22992 3482 23004
rect 6638 22992 6644 23004
rect 6696 22992 6702 23044
rect 4157 22967 4215 22973
rect 4157 22933 4169 22967
rect 4203 22964 4215 22967
rect 4706 22964 4712 22976
rect 4203 22936 4712 22964
rect 4203 22933 4215 22936
rect 4157 22927 4215 22933
rect 4706 22924 4712 22936
rect 4764 22924 4770 22976
rect 4801 22967 4859 22973
rect 4801 22933 4813 22967
rect 4847 22964 4859 22967
rect 6886 22964 6914 23072
rect 9861 23069 9873 23072
rect 9907 23069 9919 23103
rect 9861 23063 9919 23069
rect 10042 22964 10048 22976
rect 4847 22936 6914 22964
rect 10003 22936 10048 22964
rect 4847 22933 4859 22936
rect 4801 22927 4859 22933
rect 10042 22924 10048 22936
rect 10100 22924 10106 22976
rect 1104 22874 10856 22896
rect 1104 22822 4213 22874
rect 4265 22822 4277 22874
rect 4329 22822 4341 22874
rect 4393 22822 4405 22874
rect 4457 22822 4469 22874
rect 4521 22822 7477 22874
rect 7529 22822 7541 22874
rect 7593 22822 7605 22874
rect 7657 22822 7669 22874
rect 7721 22822 7733 22874
rect 7785 22822 10856 22874
rect 1104 22800 10856 22822
rect 1762 22720 1768 22772
rect 1820 22760 1826 22772
rect 2133 22763 2191 22769
rect 2133 22760 2145 22763
rect 1820 22732 2145 22760
rect 1820 22720 1826 22732
rect 2133 22729 2145 22732
rect 2179 22729 2191 22763
rect 2133 22723 2191 22729
rect 3145 22763 3203 22769
rect 3145 22729 3157 22763
rect 3191 22760 3203 22763
rect 3878 22760 3884 22772
rect 3191 22732 3884 22760
rect 3191 22729 3203 22732
rect 3145 22723 3203 22729
rect 3878 22720 3884 22732
rect 3936 22720 3942 22772
rect 4706 22720 4712 22772
rect 4764 22760 4770 22772
rect 9858 22760 9864 22772
rect 4764 22732 9864 22760
rect 4764 22720 4770 22732
rect 9858 22720 9864 22732
rect 9916 22720 9922 22772
rect 1394 22624 1400 22636
rect 1355 22596 1400 22624
rect 1394 22584 1400 22596
rect 1452 22584 1458 22636
rect 1670 22584 1676 22636
rect 1728 22624 1734 22636
rect 2041 22627 2099 22633
rect 2041 22624 2053 22627
rect 1728 22596 2053 22624
rect 1728 22584 1734 22596
rect 2041 22593 2053 22596
rect 2087 22593 2099 22627
rect 2041 22587 2099 22593
rect 2317 22627 2375 22633
rect 2317 22593 2329 22627
rect 2363 22624 2375 22627
rect 2958 22624 2964 22636
rect 2363 22596 2964 22624
rect 2363 22593 2375 22596
rect 2317 22587 2375 22593
rect 2958 22584 2964 22596
rect 3016 22584 3022 22636
rect 3237 22627 3295 22633
rect 3237 22593 3249 22627
rect 3283 22624 3295 22627
rect 4525 22627 4583 22633
rect 3283 22596 3372 22624
rect 3283 22593 3295 22596
rect 3237 22587 3295 22593
rect 1489 22559 1547 22565
rect 1489 22525 1501 22559
rect 1535 22556 1547 22559
rect 3344 22556 3372 22596
rect 4525 22593 4537 22627
rect 4571 22624 4583 22627
rect 4614 22624 4620 22636
rect 4571 22596 4620 22624
rect 4571 22593 4583 22596
rect 4525 22587 4583 22593
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 1535 22528 3372 22556
rect 1535 22525 1547 22528
rect 1489 22519 1547 22525
rect 3344 22488 3372 22528
rect 4249 22559 4307 22565
rect 4249 22525 4261 22559
rect 4295 22556 4307 22559
rect 4798 22556 4804 22568
rect 4295 22528 4804 22556
rect 4295 22525 4307 22528
rect 4249 22519 4307 22525
rect 4798 22516 4804 22528
rect 4856 22516 4862 22568
rect 4706 22488 4712 22500
rect 3344 22460 4712 22488
rect 4706 22448 4712 22460
rect 4764 22448 4770 22500
rect 1104 22330 10856 22352
rect 1104 22278 2582 22330
rect 2634 22278 2646 22330
rect 2698 22278 2710 22330
rect 2762 22278 2774 22330
rect 2826 22278 2838 22330
rect 2890 22278 5845 22330
rect 5897 22278 5909 22330
rect 5961 22278 5973 22330
rect 6025 22278 6037 22330
rect 6089 22278 6101 22330
rect 6153 22278 9109 22330
rect 9161 22278 9173 22330
rect 9225 22278 9237 22330
rect 9289 22278 9301 22330
rect 9353 22278 9365 22330
rect 9417 22278 10856 22330
rect 1104 22256 10856 22278
rect 2869 22219 2927 22225
rect 2869 22185 2881 22219
rect 2915 22216 2927 22219
rect 2958 22216 2964 22228
rect 2915 22188 2964 22216
rect 2915 22185 2927 22188
rect 2869 22179 2927 22185
rect 2958 22176 2964 22188
rect 3016 22176 3022 22228
rect 3602 22080 3608 22092
rect 1596 22052 3608 22080
rect 1596 22021 1624 22052
rect 3602 22040 3608 22052
rect 3660 22040 3666 22092
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 21981 1639 22015
rect 2038 22012 2044 22024
rect 1999 21984 2044 22012
rect 1581 21975 1639 21981
rect 2038 21972 2044 21984
rect 2096 21972 2102 22024
rect 2961 22015 3019 22021
rect 2961 21981 2973 22015
rect 3007 22012 3019 22015
rect 3050 22012 3056 22024
rect 3007 21984 3056 22012
rect 3007 21981 3019 21984
rect 2961 21975 3019 21981
rect 3050 21972 3056 21984
rect 3108 21972 3114 22024
rect 3142 21972 3148 22024
rect 3200 22012 3206 22024
rect 4065 22015 4123 22021
rect 4065 22012 4077 22015
rect 3200 21984 4077 22012
rect 3200 21972 3206 21984
rect 4065 21981 4077 21984
rect 4111 21981 4123 22015
rect 4065 21975 4123 21981
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 22012 4307 22015
rect 4614 22012 4620 22024
rect 4295 21984 4620 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 9858 22012 9864 22024
rect 9819 21984 9864 22012
rect 9858 21972 9864 21984
rect 9916 21972 9922 22024
rect 1489 21879 1547 21885
rect 1489 21845 1501 21879
rect 1535 21876 1547 21879
rect 1670 21876 1676 21888
rect 1535 21848 1676 21876
rect 1535 21845 1547 21848
rect 1489 21839 1547 21845
rect 1670 21836 1676 21848
rect 1728 21836 1734 21888
rect 2225 21879 2283 21885
rect 2225 21845 2237 21879
rect 2271 21876 2283 21879
rect 2498 21876 2504 21888
rect 2271 21848 2504 21876
rect 2271 21845 2283 21848
rect 2225 21839 2283 21845
rect 2498 21836 2504 21848
rect 2556 21836 2562 21888
rect 4157 21879 4215 21885
rect 4157 21845 4169 21879
rect 4203 21876 4215 21879
rect 9858 21876 9864 21888
rect 4203 21848 9864 21876
rect 4203 21845 4215 21848
rect 4157 21839 4215 21845
rect 9858 21836 9864 21848
rect 9916 21836 9922 21888
rect 10042 21876 10048 21888
rect 10003 21848 10048 21876
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 1104 21786 10856 21808
rect 1104 21734 4213 21786
rect 4265 21734 4277 21786
rect 4329 21734 4341 21786
rect 4393 21734 4405 21786
rect 4457 21734 4469 21786
rect 4521 21734 7477 21786
rect 7529 21734 7541 21786
rect 7593 21734 7605 21786
rect 7657 21734 7669 21786
rect 7721 21734 7733 21786
rect 7785 21734 10856 21786
rect 1104 21712 10856 21734
rect 1394 21632 1400 21684
rect 1452 21672 1458 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1452 21644 1593 21672
rect 1452 21632 1458 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 1581 21635 1639 21641
rect 1670 21564 1676 21616
rect 1728 21604 1734 21616
rect 1728 21576 4108 21604
rect 1728 21564 1734 21576
rect 1397 21539 1455 21545
rect 1397 21505 1409 21539
rect 1443 21536 1455 21539
rect 1486 21536 1492 21548
rect 1443 21508 1492 21536
rect 1443 21505 1455 21508
rect 1397 21499 1455 21505
rect 1486 21496 1492 21508
rect 1544 21496 1550 21548
rect 1578 21496 1584 21548
rect 1636 21536 1642 21548
rect 2225 21539 2283 21545
rect 2225 21536 2237 21539
rect 1636 21508 2237 21536
rect 1636 21496 1642 21508
rect 2225 21505 2237 21508
rect 2271 21505 2283 21539
rect 2866 21536 2872 21548
rect 2827 21508 2872 21536
rect 2225 21499 2283 21505
rect 2866 21496 2872 21508
rect 2924 21496 2930 21548
rect 3326 21536 3332 21548
rect 3287 21508 3332 21536
rect 3326 21496 3332 21508
rect 3384 21496 3390 21548
rect 4080 21545 4108 21576
rect 4632 21576 4936 21604
rect 4632 21548 4660 21576
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 4249 21539 4307 21545
rect 4249 21505 4261 21539
rect 4295 21536 4307 21539
rect 4614 21536 4620 21548
rect 4295 21508 4620 21536
rect 4295 21505 4307 21508
rect 4249 21499 4307 21505
rect 4614 21496 4620 21508
rect 4672 21496 4678 21548
rect 4706 21496 4712 21548
rect 4764 21536 4770 21548
rect 4908 21545 4936 21576
rect 4893 21539 4951 21545
rect 4764 21508 4809 21536
rect 4764 21496 4770 21508
rect 4893 21505 4905 21539
rect 4939 21505 4951 21539
rect 4893 21499 4951 21505
rect 4249 21403 4307 21409
rect 4249 21369 4261 21403
rect 4295 21400 4307 21403
rect 10965 21403 11023 21409
rect 10965 21400 10977 21403
rect 4295 21372 10977 21400
rect 4295 21369 4307 21372
rect 4249 21363 4307 21369
rect 10965 21369 10977 21372
rect 11011 21369 11023 21403
rect 10965 21363 11023 21369
rect 1854 21292 1860 21344
rect 1912 21332 1918 21344
rect 2041 21335 2099 21341
rect 2041 21332 2053 21335
rect 1912 21304 2053 21332
rect 1912 21292 1918 21304
rect 2041 21301 2053 21304
rect 2087 21301 2099 21335
rect 2041 21295 2099 21301
rect 2222 21292 2228 21344
rect 2280 21332 2286 21344
rect 2685 21335 2743 21341
rect 2685 21332 2697 21335
rect 2280 21304 2697 21332
rect 2280 21292 2286 21304
rect 2685 21301 2697 21304
rect 2731 21301 2743 21335
rect 2685 21295 2743 21301
rect 3513 21335 3571 21341
rect 3513 21301 3525 21335
rect 3559 21332 3571 21335
rect 3786 21332 3792 21344
rect 3559 21304 3792 21332
rect 3559 21301 3571 21304
rect 3513 21295 3571 21301
rect 3786 21292 3792 21304
rect 3844 21292 3850 21344
rect 4890 21332 4896 21344
rect 4851 21304 4896 21332
rect 4890 21292 4896 21304
rect 4948 21292 4954 21344
rect 1104 21242 10856 21264
rect 1104 21190 2582 21242
rect 2634 21190 2646 21242
rect 2698 21190 2710 21242
rect 2762 21190 2774 21242
rect 2826 21190 2838 21242
rect 2890 21190 5845 21242
rect 5897 21190 5909 21242
rect 5961 21190 5973 21242
rect 6025 21190 6037 21242
rect 6089 21190 6101 21242
rect 6153 21190 9109 21242
rect 9161 21190 9173 21242
rect 9225 21190 9237 21242
rect 9289 21190 9301 21242
rect 9353 21190 9365 21242
rect 9417 21190 10856 21242
rect 1104 21168 10856 21190
rect 4890 21088 4896 21140
rect 4948 21128 4954 21140
rect 9766 21128 9772 21140
rect 4948 21100 9772 21128
rect 4948 21088 4954 21100
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20992 4491 20995
rect 4798 20992 4804 21004
rect 4479 20964 4804 20992
rect 4479 20961 4491 20964
rect 4433 20955 4491 20961
rect 4798 20952 4804 20964
rect 4856 20952 4862 21004
rect 1397 20927 1455 20933
rect 1397 20893 1409 20927
rect 1443 20924 1455 20927
rect 1486 20924 1492 20936
rect 1443 20896 1492 20924
rect 1443 20893 1455 20896
rect 1397 20887 1455 20893
rect 1486 20884 1492 20896
rect 1544 20884 1550 20936
rect 1670 20884 1676 20936
rect 1728 20924 1734 20936
rect 2225 20927 2283 20933
rect 2225 20924 2237 20927
rect 1728 20896 2237 20924
rect 1728 20884 1734 20896
rect 2225 20893 2237 20896
rect 2271 20893 2283 20927
rect 3050 20924 3056 20936
rect 3011 20896 3056 20924
rect 2225 20887 2283 20893
rect 3050 20884 3056 20896
rect 3108 20884 3114 20936
rect 4706 20924 4712 20936
rect 4667 20896 4712 20924
rect 4706 20884 4712 20896
rect 4764 20884 4770 20936
rect 9858 20924 9864 20936
rect 9819 20896 9864 20924
rect 9858 20884 9864 20896
rect 9916 20884 9922 20936
rect 1581 20791 1639 20797
rect 1581 20757 1593 20791
rect 1627 20788 1639 20791
rect 1762 20788 1768 20800
rect 1627 20760 1768 20788
rect 1627 20757 1639 20760
rect 1581 20751 1639 20757
rect 1762 20748 1768 20760
rect 1820 20748 1826 20800
rect 2038 20788 2044 20800
rect 1999 20760 2044 20788
rect 2038 20748 2044 20760
rect 2096 20748 2102 20800
rect 2869 20791 2927 20797
rect 2869 20757 2881 20791
rect 2915 20788 2927 20791
rect 3050 20788 3056 20800
rect 2915 20760 3056 20788
rect 2915 20757 2927 20760
rect 2869 20751 2927 20757
rect 3050 20748 3056 20760
rect 3108 20748 3114 20800
rect 10042 20788 10048 20800
rect 10003 20760 10048 20788
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 1104 20698 10856 20720
rect 1104 20646 4213 20698
rect 4265 20646 4277 20698
rect 4329 20646 4341 20698
rect 4393 20646 4405 20698
rect 4457 20646 4469 20698
rect 4521 20646 7477 20698
rect 7529 20646 7541 20698
rect 7593 20646 7605 20698
rect 7657 20646 7669 20698
rect 7721 20646 7733 20698
rect 7785 20646 10856 20698
rect 1104 20624 10856 20646
rect 2133 20519 2191 20525
rect 2133 20485 2145 20519
rect 2179 20516 2191 20519
rect 4154 20516 4160 20528
rect 2179 20488 4160 20516
rect 2179 20485 2191 20488
rect 2133 20479 2191 20485
rect 4154 20476 4160 20488
rect 4212 20476 4218 20528
rect 1394 20448 1400 20460
rect 1355 20420 1400 20448
rect 1394 20408 1400 20420
rect 1452 20408 1458 20460
rect 2222 20448 2228 20460
rect 2183 20420 2228 20448
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 2498 20408 2504 20460
rect 2556 20448 2562 20460
rect 2685 20451 2743 20457
rect 2685 20448 2697 20451
rect 2556 20420 2697 20448
rect 2556 20408 2562 20420
rect 2685 20417 2697 20420
rect 2731 20417 2743 20451
rect 3510 20448 3516 20460
rect 3471 20420 3516 20448
rect 2685 20411 2743 20417
rect 3510 20408 3516 20420
rect 3568 20408 3574 20460
rect 2406 20340 2412 20392
rect 2464 20380 2470 20392
rect 7190 20380 7196 20392
rect 2464 20352 7196 20380
rect 2464 20340 2470 20352
rect 7190 20340 7196 20352
rect 7248 20340 7254 20392
rect 2777 20315 2835 20321
rect 2777 20281 2789 20315
rect 2823 20312 2835 20315
rect 4614 20312 4620 20324
rect 2823 20284 4620 20312
rect 2823 20281 2835 20284
rect 2777 20275 2835 20281
rect 4614 20272 4620 20284
rect 4672 20272 4678 20324
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 3326 20244 3332 20256
rect 3287 20216 3332 20244
rect 3326 20204 3332 20216
rect 3384 20204 3390 20256
rect 1104 20154 10856 20176
rect 1104 20102 2582 20154
rect 2634 20102 2646 20154
rect 2698 20102 2710 20154
rect 2762 20102 2774 20154
rect 2826 20102 2838 20154
rect 2890 20102 5845 20154
rect 5897 20102 5909 20154
rect 5961 20102 5973 20154
rect 6025 20102 6037 20154
rect 6089 20102 6101 20154
rect 6153 20102 9109 20154
rect 9161 20102 9173 20154
rect 9225 20102 9237 20154
rect 9289 20102 9301 20154
rect 9353 20102 9365 20154
rect 9417 20102 10856 20154
rect 1104 20080 10856 20102
rect 7098 20040 7104 20052
rect 2424 20012 7104 20040
rect 2424 19981 2452 20012
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 2409 19975 2467 19981
rect 2409 19941 2421 19975
rect 2455 19941 2467 19975
rect 2409 19935 2467 19941
rect 2958 19932 2964 19984
rect 3016 19972 3022 19984
rect 7006 19972 7012 19984
rect 3016 19944 7012 19972
rect 3016 19932 3022 19944
rect 7006 19932 7012 19944
rect 7064 19932 7070 19984
rect 750 19864 756 19916
rect 808 19904 814 19916
rect 2130 19904 2136 19916
rect 808 19876 2136 19904
rect 808 19864 814 19876
rect 2130 19864 2136 19876
rect 2188 19864 2194 19916
rect 3050 19904 3056 19916
rect 2516 19876 3056 19904
rect 2516 19848 2544 19876
rect 3050 19864 3056 19876
rect 3108 19864 3114 19916
rect 3510 19864 3516 19916
rect 3568 19904 3574 19916
rect 5166 19904 5172 19916
rect 3568 19876 5172 19904
rect 3568 19864 3574 19876
rect 5166 19864 5172 19876
rect 5224 19864 5230 19916
rect 1854 19836 1860 19848
rect 1815 19808 1860 19836
rect 1854 19796 1860 19808
rect 1912 19796 1918 19848
rect 2498 19836 2504 19848
rect 2411 19808 2504 19836
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19836 2743 19839
rect 3142 19836 3148 19848
rect 2731 19808 3148 19836
rect 2731 19805 2743 19808
rect 2685 19799 2743 19805
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 3786 19836 3792 19848
rect 3747 19808 3792 19836
rect 3786 19796 3792 19808
rect 3844 19796 3850 19848
rect 9766 19796 9772 19848
rect 9824 19836 9830 19848
rect 9861 19839 9919 19845
rect 9861 19836 9873 19839
rect 9824 19808 9873 19836
rect 9824 19796 9830 19808
rect 9861 19805 9873 19808
rect 9907 19805 9919 19839
rect 9861 19799 9919 19805
rect 1765 19771 1823 19777
rect 1765 19737 1777 19771
rect 1811 19768 1823 19771
rect 4982 19768 4988 19780
rect 1811 19740 4988 19768
rect 1811 19737 1823 19740
rect 1765 19731 1823 19737
rect 1872 19712 1900 19740
rect 4982 19728 4988 19740
rect 5040 19728 5046 19780
rect 1854 19660 1860 19712
rect 1912 19660 1918 19712
rect 3050 19660 3056 19712
rect 3108 19700 3114 19712
rect 3881 19703 3939 19709
rect 3881 19700 3893 19703
rect 3108 19672 3893 19700
rect 3108 19660 3114 19672
rect 3881 19669 3893 19672
rect 3927 19669 3939 19703
rect 10042 19700 10048 19712
rect 10003 19672 10048 19700
rect 3881 19663 3939 19669
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 1104 19610 10856 19632
rect 1104 19558 4213 19610
rect 4265 19558 4277 19610
rect 4329 19558 4341 19610
rect 4393 19558 4405 19610
rect 4457 19558 4469 19610
rect 4521 19558 7477 19610
rect 7529 19558 7541 19610
rect 7593 19558 7605 19610
rect 7657 19558 7669 19610
rect 7721 19558 7733 19610
rect 7785 19558 10856 19610
rect 1104 19536 10856 19558
rect 1765 19499 1823 19505
rect 1765 19465 1777 19499
rect 1811 19496 1823 19499
rect 2406 19496 2412 19508
rect 1811 19468 2412 19496
rect 1811 19465 1823 19468
rect 1765 19459 1823 19465
rect 2406 19456 2412 19468
rect 2464 19456 2470 19508
rect 2958 19496 2964 19508
rect 2919 19468 2964 19496
rect 2958 19456 2964 19468
rect 3016 19456 3022 19508
rect 3789 19499 3847 19505
rect 3789 19465 3801 19499
rect 3835 19496 3847 19499
rect 3970 19496 3976 19508
rect 3835 19468 3976 19496
rect 3835 19465 3847 19468
rect 3789 19459 3847 19465
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 4614 19428 4620 19440
rect 1688 19400 2544 19428
rect 1688 19369 1716 19400
rect 2516 19372 2544 19400
rect 3068 19400 4620 19428
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19329 1731 19363
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1673 19323 1731 19329
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 2498 19360 2504 19372
rect 2459 19332 2504 19360
rect 2498 19320 2504 19332
rect 2556 19360 2562 19372
rect 3068 19369 3096 19400
rect 4614 19388 4620 19400
rect 4672 19388 4678 19440
rect 3053 19363 3111 19369
rect 2556 19332 3004 19360
rect 2556 19320 2562 19332
rect 2976 19292 3004 19332
rect 3053 19329 3065 19363
rect 3099 19329 3111 19363
rect 3605 19363 3663 19369
rect 3605 19360 3617 19363
rect 3053 19323 3111 19329
rect 3160 19332 3617 19360
rect 3160 19292 3188 19332
rect 3605 19329 3617 19332
rect 3651 19329 3663 19363
rect 3605 19323 3663 19329
rect 3881 19363 3939 19369
rect 3881 19329 3893 19363
rect 3927 19360 3939 19363
rect 4062 19360 4068 19372
rect 3927 19332 4068 19360
rect 3927 19329 3939 19332
rect 3881 19323 3939 19329
rect 4062 19320 4068 19332
rect 4120 19360 4126 19372
rect 4798 19360 4804 19372
rect 4120 19332 4804 19360
rect 4120 19320 4126 19332
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 2976 19264 3188 19292
rect 2958 19184 2964 19236
rect 3016 19224 3022 19236
rect 3418 19224 3424 19236
rect 3016 19196 3424 19224
rect 3016 19184 3022 19196
rect 3418 19184 3424 19196
rect 3476 19184 3482 19236
rect 1104 19066 10856 19088
rect 1104 19014 2582 19066
rect 2634 19014 2646 19066
rect 2698 19014 2710 19066
rect 2762 19014 2774 19066
rect 2826 19014 2838 19066
rect 2890 19014 5845 19066
rect 5897 19014 5909 19066
rect 5961 19014 5973 19066
rect 6025 19014 6037 19066
rect 6089 19014 6101 19066
rect 6153 19014 9109 19066
rect 9161 19014 9173 19066
rect 9225 19014 9237 19066
rect 9289 19014 9301 19066
rect 9353 19014 9365 19066
rect 9417 19014 10856 19066
rect 1104 18992 10856 19014
rect 1765 18955 1823 18961
rect 1765 18921 1777 18955
rect 1811 18952 1823 18955
rect 3510 18952 3516 18964
rect 1811 18924 3516 18952
rect 1811 18921 1823 18924
rect 1765 18915 1823 18921
rect 3510 18912 3516 18924
rect 3568 18912 3574 18964
rect 1857 18751 1915 18757
rect 1857 18717 1869 18751
rect 1903 18748 1915 18751
rect 2038 18748 2044 18760
rect 1903 18720 2044 18748
rect 1903 18717 1915 18720
rect 1857 18711 1915 18717
rect 2038 18708 2044 18720
rect 2096 18708 2102 18760
rect 2498 18748 2504 18760
rect 2459 18720 2504 18748
rect 2498 18708 2504 18720
rect 2556 18708 2562 18760
rect 3050 18748 3056 18760
rect 3011 18720 3056 18748
rect 3050 18708 3056 18720
rect 3108 18708 3114 18760
rect 3970 18748 3976 18760
rect 3931 18720 3976 18748
rect 3970 18708 3976 18720
rect 4028 18708 4034 18760
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18748 9919 18751
rect 10965 18751 11023 18757
rect 10965 18748 10977 18751
rect 9907 18720 10977 18748
rect 9907 18717 9919 18720
rect 9861 18711 9919 18717
rect 10965 18717 10977 18720
rect 11011 18717 11023 18751
rect 10965 18711 11023 18717
rect 7834 18680 7840 18692
rect 2976 18652 7840 18680
rect 2976 18621 3004 18652
rect 7834 18640 7840 18652
rect 7892 18640 7898 18692
rect 2961 18615 3019 18621
rect 2961 18581 2973 18615
rect 3007 18581 3019 18615
rect 3786 18612 3792 18624
rect 3747 18584 3792 18612
rect 2961 18575 3019 18581
rect 3786 18572 3792 18584
rect 3844 18572 3850 18624
rect 10042 18612 10048 18624
rect 10003 18584 10048 18612
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 1104 18522 10856 18544
rect 1104 18470 4213 18522
rect 4265 18470 4277 18522
rect 4329 18470 4341 18522
rect 4393 18470 4405 18522
rect 4457 18470 4469 18522
rect 4521 18470 7477 18522
rect 7529 18470 7541 18522
rect 7593 18470 7605 18522
rect 7657 18470 7669 18522
rect 7721 18470 7733 18522
rect 7785 18470 10856 18522
rect 1104 18448 10856 18470
rect 2130 18408 2136 18420
rect 2091 18380 2136 18408
rect 2130 18368 2136 18380
rect 2188 18368 2194 18420
rect 4614 18340 4620 18352
rect 4356 18312 4620 18340
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 1762 18232 1768 18284
rect 1820 18272 1826 18284
rect 2041 18275 2099 18281
rect 2041 18272 2053 18275
rect 1820 18244 2053 18272
rect 1820 18232 1826 18244
rect 2041 18241 2053 18244
rect 2087 18241 2099 18275
rect 2041 18235 2099 18241
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18272 2927 18275
rect 3326 18272 3332 18284
rect 2915 18244 3332 18272
rect 2915 18241 2927 18244
rect 2869 18235 2927 18241
rect 3326 18232 3332 18244
rect 3384 18232 3390 18284
rect 3510 18272 3516 18284
rect 3471 18244 3516 18272
rect 3510 18232 3516 18244
rect 3568 18232 3574 18284
rect 4356 18281 4384 18312
rect 4614 18300 4620 18312
rect 4672 18300 4678 18352
rect 4724 18312 5212 18340
rect 4724 18284 4752 18312
rect 4341 18275 4399 18281
rect 4341 18241 4353 18275
rect 4387 18241 4399 18275
rect 4341 18235 4399 18241
rect 4525 18275 4583 18281
rect 4525 18241 4537 18275
rect 4571 18272 4583 18275
rect 4706 18272 4712 18284
rect 4571 18244 4712 18272
rect 4571 18241 4583 18244
rect 4525 18235 4583 18241
rect 4706 18232 4712 18244
rect 4764 18232 4770 18284
rect 5184 18281 5212 18312
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18241 5043 18275
rect 4985 18235 5043 18241
rect 5169 18275 5227 18281
rect 5169 18241 5181 18275
rect 5215 18241 5227 18275
rect 5169 18235 5227 18241
rect 3050 18164 3056 18216
rect 3108 18204 3114 18216
rect 5000 18204 5028 18235
rect 3108 18176 5028 18204
rect 3108 18164 3114 18176
rect 842 18096 848 18148
rect 900 18136 906 18148
rect 2038 18136 2044 18148
rect 900 18108 2044 18136
rect 900 18096 906 18108
rect 2038 18096 2044 18108
rect 2096 18096 2102 18148
rect 2777 18139 2835 18145
rect 2777 18105 2789 18139
rect 2823 18136 2835 18139
rect 3142 18136 3148 18148
rect 2823 18108 3148 18136
rect 2823 18105 2835 18108
rect 2777 18099 2835 18105
rect 3142 18096 3148 18108
rect 3200 18136 3206 18148
rect 4338 18136 4344 18148
rect 3200 18108 4344 18136
rect 3200 18096 3206 18108
rect 4338 18096 4344 18108
rect 4396 18096 4402 18148
rect 4525 18139 4583 18145
rect 4525 18105 4537 18139
rect 4571 18136 4583 18139
rect 9766 18136 9772 18148
rect 4571 18108 9772 18136
rect 4571 18105 4583 18108
rect 4525 18099 4583 18105
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 1486 18028 1492 18080
rect 1544 18068 1550 18080
rect 1581 18071 1639 18077
rect 1581 18068 1593 18071
rect 1544 18040 1593 18068
rect 1544 18028 1550 18040
rect 1581 18037 1593 18040
rect 1627 18037 1639 18071
rect 1581 18031 1639 18037
rect 2130 18028 2136 18080
rect 2188 18068 2194 18080
rect 3050 18068 3056 18080
rect 2188 18040 3056 18068
rect 2188 18028 2194 18040
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 3326 18068 3332 18080
rect 3287 18040 3332 18068
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 5169 18071 5227 18077
rect 5169 18037 5181 18071
rect 5215 18068 5227 18071
rect 9858 18068 9864 18080
rect 5215 18040 9864 18068
rect 5215 18037 5227 18040
rect 5169 18031 5227 18037
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 1104 17978 10856 18000
rect 1104 17926 2582 17978
rect 2634 17926 2646 17978
rect 2698 17926 2710 17978
rect 2762 17926 2774 17978
rect 2826 17926 2838 17978
rect 2890 17926 5845 17978
rect 5897 17926 5909 17978
rect 5961 17926 5973 17978
rect 6025 17926 6037 17978
rect 6089 17926 6101 17978
rect 6153 17926 9109 17978
rect 9161 17926 9173 17978
rect 9225 17926 9237 17978
rect 9289 17926 9301 17978
rect 9353 17926 9365 17978
rect 9417 17926 10856 17978
rect 1104 17904 10856 17926
rect 2133 17867 2191 17873
rect 2133 17833 2145 17867
rect 2179 17864 2191 17867
rect 3970 17864 3976 17876
rect 2179 17836 3976 17864
rect 2179 17833 2191 17836
rect 2133 17827 2191 17833
rect 3970 17824 3976 17836
rect 4028 17864 4034 17876
rect 6454 17864 6460 17876
rect 4028 17836 6460 17864
rect 4028 17824 4034 17836
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 934 17620 940 17672
rect 992 17660 998 17672
rect 1397 17663 1455 17669
rect 1397 17660 1409 17663
rect 992 17632 1409 17660
rect 992 17620 998 17632
rect 1397 17629 1409 17632
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 1578 17620 1584 17672
rect 1636 17660 1642 17672
rect 2041 17663 2099 17669
rect 2041 17660 2053 17663
rect 1636 17632 2053 17660
rect 1636 17620 1642 17632
rect 2041 17629 2053 17632
rect 2087 17629 2099 17663
rect 2866 17660 2872 17672
rect 2827 17632 2872 17660
rect 2041 17623 2099 17629
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 4338 17660 4344 17672
rect 4299 17632 4344 17660
rect 4338 17620 4344 17632
rect 4396 17620 4402 17672
rect 4525 17663 4583 17669
rect 4525 17629 4537 17663
rect 4571 17660 4583 17663
rect 4706 17660 4712 17672
rect 4571 17632 4712 17660
rect 4571 17629 4583 17632
rect 4525 17623 4583 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 4982 17660 4988 17672
rect 4943 17632 4988 17660
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5169 17663 5227 17669
rect 5169 17629 5181 17663
rect 5215 17629 5227 17663
rect 9858 17660 9864 17672
rect 9819 17632 9864 17660
rect 5169 17623 5227 17629
rect 4724 17592 4752 17620
rect 5184 17592 5212 17623
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 10965 17595 11023 17601
rect 10965 17592 10977 17595
rect 4724 17564 5212 17592
rect 6886 17564 10977 17592
rect 1578 17524 1584 17536
rect 1539 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 2222 17484 2228 17536
rect 2280 17524 2286 17536
rect 2685 17527 2743 17533
rect 2685 17524 2697 17527
rect 2280 17496 2697 17524
rect 2280 17484 2286 17496
rect 2685 17493 2697 17496
rect 2731 17493 2743 17527
rect 2685 17487 2743 17493
rect 4433 17527 4491 17533
rect 4433 17493 4445 17527
rect 4479 17524 4491 17527
rect 4982 17524 4988 17536
rect 4479 17496 4988 17524
rect 4479 17493 4491 17496
rect 4433 17487 4491 17493
rect 4982 17484 4988 17496
rect 5040 17484 5046 17536
rect 5077 17527 5135 17533
rect 5077 17493 5089 17527
rect 5123 17524 5135 17527
rect 6886 17524 6914 17564
rect 10965 17561 10977 17564
rect 11011 17561 11023 17595
rect 10965 17555 11023 17561
rect 10042 17524 10048 17536
rect 5123 17496 6914 17524
rect 10003 17496 10048 17524
rect 5123 17493 5135 17496
rect 5077 17487 5135 17493
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 1104 17434 10856 17456
rect 1104 17382 4213 17434
rect 4265 17382 4277 17434
rect 4329 17382 4341 17434
rect 4393 17382 4405 17434
rect 4457 17382 4469 17434
rect 4521 17382 7477 17434
rect 7529 17382 7541 17434
rect 7593 17382 7605 17434
rect 7657 17382 7669 17434
rect 7721 17382 7733 17434
rect 7785 17382 10856 17434
rect 1104 17360 10856 17382
rect 2038 17280 2044 17332
rect 2096 17320 2102 17332
rect 2133 17323 2191 17329
rect 2133 17320 2145 17323
rect 2096 17292 2145 17320
rect 2096 17280 2102 17292
rect 2133 17289 2145 17292
rect 2179 17320 2191 17323
rect 3694 17320 3700 17332
rect 2179 17292 3700 17320
rect 2179 17289 2191 17292
rect 2133 17283 2191 17289
rect 3694 17280 3700 17292
rect 3752 17280 3758 17332
rect 4982 17280 4988 17332
rect 5040 17320 5046 17332
rect 11057 17323 11115 17329
rect 11057 17320 11069 17323
rect 5040 17292 11069 17320
rect 5040 17280 5046 17292
rect 11057 17289 11069 17292
rect 11103 17289 11115 17323
rect 11057 17283 11115 17289
rect 4798 17252 4804 17264
rect 4356 17224 4804 17252
rect 1394 17184 1400 17196
rect 1355 17156 1400 17184
rect 1394 17144 1400 17156
rect 1452 17144 1458 17196
rect 2225 17187 2283 17193
rect 2225 17153 2237 17187
rect 2271 17184 2283 17187
rect 3786 17184 3792 17196
rect 2271 17156 3792 17184
rect 2271 17153 2283 17156
rect 2225 17147 2283 17153
rect 3786 17144 3792 17156
rect 3844 17144 3850 17196
rect 4356 17193 4384 17224
rect 4798 17212 4804 17224
rect 4856 17212 4862 17264
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17153 4399 17187
rect 4341 17147 4399 17153
rect 4525 17187 4583 17193
rect 4525 17153 4537 17187
rect 4571 17184 4583 17187
rect 4706 17184 4712 17196
rect 4571 17156 4712 17184
rect 4571 17153 4583 17156
rect 4525 17147 4583 17153
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 1581 16983 1639 16989
rect 1581 16949 1593 16983
rect 1627 16980 1639 16983
rect 1670 16980 1676 16992
rect 1627 16952 1676 16980
rect 1627 16949 1639 16952
rect 1581 16943 1639 16949
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 4525 16983 4583 16989
rect 4525 16949 4537 16983
rect 4571 16980 4583 16983
rect 9858 16980 9864 16992
rect 4571 16952 9864 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 1104 16890 10856 16912
rect 1104 16838 2582 16890
rect 2634 16838 2646 16890
rect 2698 16838 2710 16890
rect 2762 16838 2774 16890
rect 2826 16838 2838 16890
rect 2890 16838 5845 16890
rect 5897 16838 5909 16890
rect 5961 16838 5973 16890
rect 6025 16838 6037 16890
rect 6089 16838 6101 16890
rect 6153 16838 9109 16890
rect 9161 16838 9173 16890
rect 9225 16838 9237 16890
rect 9289 16838 9301 16890
rect 9353 16838 9365 16890
rect 9417 16838 10856 16890
rect 1104 16816 10856 16838
rect 1949 16779 2007 16785
rect 1949 16745 1961 16779
rect 1995 16776 2007 16779
rect 2222 16776 2228 16788
rect 1995 16748 2228 16776
rect 1995 16745 2007 16748
rect 1949 16739 2007 16745
rect 2222 16736 2228 16748
rect 2280 16736 2286 16788
rect 1486 16640 1492 16652
rect 1447 16612 1492 16640
rect 1486 16600 1492 16612
rect 1544 16600 1550 16652
rect 1578 16572 1584 16584
rect 1539 16544 1584 16572
rect 1578 16532 1584 16544
rect 1636 16532 1642 16584
rect 1949 16575 2007 16581
rect 1949 16541 1961 16575
rect 1995 16572 2007 16575
rect 3326 16572 3332 16584
rect 1995 16544 3332 16572
rect 1995 16541 2007 16544
rect 1949 16535 2007 16541
rect 3326 16532 3332 16544
rect 3384 16532 3390 16584
rect 9766 16532 9772 16584
rect 9824 16572 9830 16584
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 9824 16544 9873 16572
rect 9824 16532 9830 16544
rect 9861 16541 9873 16544
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 2130 16436 2136 16448
rect 2091 16408 2136 16436
rect 2130 16396 2136 16408
rect 2188 16396 2194 16448
rect 10042 16436 10048 16448
rect 10003 16408 10048 16436
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 1104 16346 10856 16368
rect 1104 16294 4213 16346
rect 4265 16294 4277 16346
rect 4329 16294 4341 16346
rect 4393 16294 4405 16346
rect 4457 16294 4469 16346
rect 4521 16294 7477 16346
rect 7529 16294 7541 16346
rect 7593 16294 7605 16346
rect 7657 16294 7669 16346
rect 7721 16294 7733 16346
rect 7785 16294 10856 16346
rect 1104 16272 10856 16294
rect 1397 16099 1455 16105
rect 1397 16065 1409 16099
rect 1443 16096 1455 16099
rect 1486 16096 1492 16108
rect 1443 16068 1492 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1486 16056 1492 16068
rect 1544 16056 1550 16108
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 1946 15960 1952 15972
rect 1627 15932 1952 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 1946 15920 1952 15932
rect 2004 15920 2010 15972
rect 1854 15852 1860 15904
rect 1912 15892 1918 15904
rect 2041 15895 2099 15901
rect 2041 15892 2053 15895
rect 1912 15864 2053 15892
rect 1912 15852 1918 15864
rect 2041 15861 2053 15864
rect 2087 15861 2099 15895
rect 2041 15855 2099 15861
rect 1104 15802 10856 15824
rect 1104 15750 2582 15802
rect 2634 15750 2646 15802
rect 2698 15750 2710 15802
rect 2762 15750 2774 15802
rect 2826 15750 2838 15802
rect 2890 15750 5845 15802
rect 5897 15750 5909 15802
rect 5961 15750 5973 15802
rect 6025 15750 6037 15802
rect 6089 15750 6101 15802
rect 6153 15750 9109 15802
rect 9161 15750 9173 15802
rect 9225 15750 9237 15802
rect 9289 15750 9301 15802
rect 9353 15750 9365 15802
rect 9417 15750 10856 15802
rect 1104 15728 10856 15750
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 2222 15484 2228 15496
rect 2183 15456 2228 15484
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 9858 15484 9864 15496
rect 9819 15456 9864 15484
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 2038 15348 2044 15360
rect 1999 15320 2044 15348
rect 2038 15308 2044 15320
rect 2096 15308 2102 15360
rect 10042 15348 10048 15360
rect 10003 15320 10048 15348
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 1104 15258 10856 15280
rect 1104 15206 4213 15258
rect 4265 15206 4277 15258
rect 4329 15206 4341 15258
rect 4393 15206 4405 15258
rect 4457 15206 4469 15258
rect 4521 15206 7477 15258
rect 7529 15206 7541 15258
rect 7593 15206 7605 15258
rect 7657 15206 7669 15258
rect 7721 15206 7733 15258
rect 7785 15206 10856 15258
rect 1104 15184 10856 15206
rect 1581 15079 1639 15085
rect 1581 15045 1593 15079
rect 1627 15076 1639 15079
rect 2038 15076 2044 15088
rect 1627 15048 2044 15076
rect 1627 15045 1639 15048
rect 1581 15039 1639 15045
rect 2038 15036 2044 15048
rect 2096 15036 2102 15088
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 15008 1455 15011
rect 1670 15008 1676 15020
rect 1443 14980 1676 15008
rect 1443 14977 1455 14980
rect 1397 14971 1455 14977
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 1762 14804 1768 14816
rect 1723 14776 1768 14804
rect 1762 14764 1768 14776
rect 1820 14764 1826 14816
rect 1104 14714 10856 14736
rect 1104 14662 2582 14714
rect 2634 14662 2646 14714
rect 2698 14662 2710 14714
rect 2762 14662 2774 14714
rect 2826 14662 2838 14714
rect 2890 14662 5845 14714
rect 5897 14662 5909 14714
rect 5961 14662 5973 14714
rect 6025 14662 6037 14714
rect 6089 14662 6101 14714
rect 6153 14662 9109 14714
rect 9161 14662 9173 14714
rect 9225 14662 9237 14714
rect 9289 14662 9301 14714
rect 9353 14662 9365 14714
rect 9417 14662 10856 14714
rect 1104 14640 10856 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 1397 14535 1455 14541
rect 1397 14501 1409 14535
rect 1443 14532 1455 14535
rect 2406 14532 2412 14544
rect 1443 14504 2412 14532
rect 1443 14501 1455 14504
rect 1397 14495 1455 14501
rect 2406 14492 2412 14504
rect 2464 14492 2470 14544
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14365 1639 14399
rect 1581 14359 1639 14365
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14396 1915 14399
rect 2130 14396 2136 14408
rect 1903 14368 2136 14396
rect 1903 14365 1915 14368
rect 1857 14359 1915 14365
rect 1596 14328 1624 14359
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 2314 14396 2320 14408
rect 2275 14368 2320 14396
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14396 9919 14399
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 9907 14368 10977 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 10965 14365 10977 14368
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 1946 14328 1952 14340
rect 1596 14300 1952 14328
rect 1946 14288 1952 14300
rect 2004 14328 2010 14340
rect 2004 14300 2176 14328
rect 2004 14288 2010 14300
rect 2148 14272 2176 14300
rect 2130 14220 2136 14272
rect 2188 14220 2194 14272
rect 2498 14260 2504 14272
rect 2459 14232 2504 14260
rect 2498 14220 2504 14232
rect 2556 14220 2562 14272
rect 10042 14260 10048 14272
rect 10003 14232 10048 14260
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 1104 14170 10856 14192
rect 1104 14118 4213 14170
rect 4265 14118 4277 14170
rect 4329 14118 4341 14170
rect 4393 14118 4405 14170
rect 4457 14118 4469 14170
rect 4521 14118 7477 14170
rect 7529 14118 7541 14170
rect 7593 14118 7605 14170
rect 7657 14118 7669 14170
rect 7721 14118 7733 14170
rect 7785 14118 10856 14170
rect 1104 14096 10856 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1670 14056 1676 14068
rect 1627 14028 1676 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 1946 14016 1952 14068
rect 2004 14056 2010 14068
rect 2041 14059 2099 14065
rect 2041 14056 2053 14059
rect 2004 14028 2053 14056
rect 2004 14016 2010 14028
rect 2041 14025 2053 14028
rect 2087 14025 2099 14059
rect 2041 14019 2099 14025
rect 1394 13920 1400 13932
rect 1355 13892 1400 13920
rect 1394 13880 1400 13892
rect 1452 13880 1458 13932
rect 2222 13920 2228 13932
rect 2183 13892 2228 13920
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 1104 13626 10856 13648
rect 1104 13574 2582 13626
rect 2634 13574 2646 13626
rect 2698 13574 2710 13626
rect 2762 13574 2774 13626
rect 2826 13574 2838 13626
rect 2890 13574 5845 13626
rect 5897 13574 5909 13626
rect 5961 13574 5973 13626
rect 6025 13574 6037 13626
rect 6089 13574 6101 13626
rect 6153 13574 9109 13626
rect 9161 13574 9173 13626
rect 9225 13574 9237 13626
rect 9289 13574 9301 13626
rect 9353 13574 9365 13626
rect 9417 13574 10856 13626
rect 1104 13552 10856 13574
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 1486 13308 1492 13320
rect 1443 13280 1492 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 1486 13268 1492 13280
rect 1544 13268 1550 13320
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 1762 13172 1768 13184
rect 1627 13144 1768 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 1104 13082 10856 13104
rect 1104 13030 4213 13082
rect 4265 13030 4277 13082
rect 4329 13030 4341 13082
rect 4393 13030 4405 13082
rect 4457 13030 4469 13082
rect 4521 13030 7477 13082
rect 7529 13030 7541 13082
rect 7593 13030 7605 13082
rect 7657 13030 7669 13082
rect 7721 13030 7733 13082
rect 7785 13030 10856 13082
rect 1104 13008 10856 13030
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 2222 12832 2228 12844
rect 2183 12804 2228 12832
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12832 9919 12835
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 9907 12804 11069 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 11057 12801 11069 12804
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 10042 12696 10048 12708
rect 10003 12668 10048 12696
rect 10042 12656 10048 12668
rect 10100 12656 10106 12708
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 1104 12538 10856 12560
rect 1104 12486 2582 12538
rect 2634 12486 2646 12538
rect 2698 12486 2710 12538
rect 2762 12486 2774 12538
rect 2826 12486 2838 12538
rect 2890 12486 5845 12538
rect 5897 12486 5909 12538
rect 5961 12486 5973 12538
rect 6025 12486 6037 12538
rect 6089 12486 6101 12538
rect 6153 12486 9109 12538
rect 9161 12486 9173 12538
rect 9225 12486 9237 12538
rect 9289 12486 9301 12538
rect 9353 12486 9365 12538
rect 9417 12486 10856 12538
rect 1104 12464 10856 12486
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 1854 12180 1860 12232
rect 1912 12220 1918 12232
rect 2225 12223 2283 12229
rect 2225 12220 2237 12223
rect 1912 12192 2237 12220
rect 1912 12180 1918 12192
rect 2225 12189 2237 12192
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 1397 12155 1455 12161
rect 1397 12121 1409 12155
rect 1443 12152 1455 12155
rect 1670 12152 1676 12164
rect 1443 12124 1676 12152
rect 1443 12121 1455 12124
rect 1397 12115 1455 12121
rect 1670 12112 1676 12124
rect 1728 12112 1734 12164
rect 1578 12044 1584 12096
rect 1636 12084 1642 12096
rect 1765 12087 1823 12093
rect 1765 12084 1777 12087
rect 1636 12056 1777 12084
rect 1636 12044 1642 12056
rect 1765 12053 1777 12056
rect 1811 12053 1823 12087
rect 1765 12047 1823 12053
rect 1854 12044 1860 12096
rect 1912 12084 1918 12096
rect 2317 12087 2375 12093
rect 2317 12084 2329 12087
rect 1912 12056 2329 12084
rect 1912 12044 1918 12056
rect 2317 12053 2329 12056
rect 2363 12053 2375 12087
rect 2317 12047 2375 12053
rect 1104 11994 10856 12016
rect 1104 11942 4213 11994
rect 4265 11942 4277 11994
rect 4329 11942 4341 11994
rect 4393 11942 4405 11994
rect 4457 11942 4469 11994
rect 4521 11942 7477 11994
rect 7529 11942 7541 11994
rect 7593 11942 7605 11994
rect 7657 11942 7669 11994
rect 7721 11942 7733 11994
rect 7785 11942 10856 11994
rect 1104 11920 10856 11942
rect 1857 11883 1915 11889
rect 1857 11849 1869 11883
rect 1903 11849 1915 11883
rect 1857 11843 1915 11849
rect 1872 11812 1900 11843
rect 2406 11812 2412 11824
rect 1872 11784 2412 11812
rect 2406 11772 2412 11784
rect 2464 11812 2470 11824
rect 2685 11815 2743 11821
rect 2685 11812 2697 11815
rect 2464 11784 2697 11812
rect 2464 11772 2470 11784
rect 2685 11781 2697 11784
rect 2731 11781 2743 11815
rect 2685 11775 2743 11781
rect 1397 11747 1455 11753
rect 1397 11713 1409 11747
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 1854 11744 1860 11756
rect 1719 11716 1860 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 1412 11608 1440 11707
rect 1854 11704 1860 11716
rect 1912 11704 1918 11756
rect 2130 11704 2136 11756
rect 2188 11744 2194 11756
rect 2317 11747 2375 11753
rect 2317 11744 2329 11747
rect 2188 11716 2329 11744
rect 2188 11704 2194 11716
rect 2317 11713 2329 11716
rect 2363 11713 2375 11747
rect 2317 11707 2375 11713
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3476 11716 3985 11744
rect 3476 11704 3482 11716
rect 3973 11713 3985 11716
rect 4019 11713 4031 11747
rect 4154 11744 4160 11756
rect 4115 11716 4160 11744
rect 3973 11707 4031 11713
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 9861 11747 9919 11753
rect 9861 11713 9873 11747
rect 9907 11713 9919 11747
rect 9861 11707 9919 11713
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11676 1639 11679
rect 2038 11676 2044 11688
rect 1627 11648 2044 11676
rect 1627 11645 1639 11648
rect 1581 11639 1639 11645
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 2409 11679 2467 11685
rect 2409 11676 2421 11679
rect 2148 11648 2421 11676
rect 1946 11608 1952 11620
rect 1412 11580 1952 11608
rect 1946 11568 1952 11580
rect 2004 11568 2010 11620
rect 1673 11543 1731 11549
rect 1673 11509 1685 11543
rect 1719 11540 1731 11543
rect 1762 11540 1768 11552
rect 1719 11512 1768 11540
rect 1719 11509 1731 11512
rect 1673 11503 1731 11509
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 2038 11500 2044 11552
rect 2096 11540 2102 11552
rect 2148 11540 2176 11648
rect 2409 11645 2421 11648
rect 2455 11676 2467 11679
rect 2498 11676 2504 11688
rect 2455 11648 2504 11676
rect 2455 11645 2467 11648
rect 2409 11639 2467 11645
rect 2498 11636 2504 11648
rect 2556 11636 2562 11688
rect 9876 11676 9904 11707
rect 4172 11648 9904 11676
rect 4172 11617 4200 11648
rect 2685 11611 2743 11617
rect 2685 11608 2697 11611
rect 2332 11580 2697 11608
rect 2332 11552 2360 11580
rect 2685 11577 2697 11580
rect 2731 11577 2743 11611
rect 2685 11571 2743 11577
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11577 4215 11611
rect 10042 11608 10048 11620
rect 10003 11580 10048 11608
rect 4157 11571 4215 11577
rect 10042 11568 10048 11580
rect 10100 11568 10106 11620
rect 2096 11512 2176 11540
rect 2096 11500 2102 11512
rect 2314 11500 2320 11552
rect 2372 11500 2378 11552
rect 2498 11500 2504 11552
rect 2556 11540 2562 11552
rect 2556 11512 2601 11540
rect 2556 11500 2562 11512
rect 1104 11450 10856 11472
rect 1104 11398 2582 11450
rect 2634 11398 2646 11450
rect 2698 11398 2710 11450
rect 2762 11398 2774 11450
rect 2826 11398 2838 11450
rect 2890 11398 5845 11450
rect 5897 11398 5909 11450
rect 5961 11398 5973 11450
rect 6025 11398 6037 11450
rect 6089 11398 6101 11450
rect 6153 11398 9109 11450
rect 9161 11398 9173 11450
rect 9225 11398 9237 11450
rect 9289 11398 9301 11450
rect 9353 11398 9365 11450
rect 9417 11398 10856 11450
rect 1104 11376 10856 11398
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 2498 11336 2504 11348
rect 1728 11308 2504 11336
rect 1728 11296 1734 11308
rect 2498 11296 2504 11308
rect 2556 11296 2562 11348
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 2958 11200 2964 11212
rect 2731 11172 2964 11200
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 5258 11200 5264 11212
rect 3936 11172 5264 11200
rect 3936 11160 3942 11172
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2130 11132 2136 11144
rect 2091 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2280 11104 2325 11132
rect 2280 11092 2286 11104
rect 2406 11092 2412 11144
rect 2464 11132 2470 11144
rect 2464 11104 2509 11132
rect 2464 11092 2470 11104
rect 3050 11092 3056 11144
rect 3108 11132 3114 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3108 11104 3985 11132
rect 3108 11092 3114 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4614 11132 4620 11144
rect 4212 11104 4620 11132
rect 4212 11092 4218 11104
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 106 11024 112 11076
rect 164 11064 170 11076
rect 2958 11064 2964 11076
rect 164 11036 2964 11064
rect 164 11024 170 11036
rect 2958 11024 2964 11036
rect 3016 11024 3022 11076
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11064 4123 11067
rect 9858 11064 9864 11076
rect 4111 11036 9864 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 1578 10996 1584 11008
rect 1539 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 1104 10906 10856 10928
rect 1104 10854 4213 10906
rect 4265 10854 4277 10906
rect 4329 10854 4341 10906
rect 4393 10854 4405 10906
rect 4457 10854 4469 10906
rect 4521 10854 7477 10906
rect 7529 10854 7541 10906
rect 7593 10854 7605 10906
rect 7657 10854 7669 10906
rect 7721 10854 7733 10906
rect 7785 10854 10856 10906
rect 1104 10832 10856 10854
rect 2685 10795 2743 10801
rect 2685 10761 2697 10795
rect 2731 10792 2743 10795
rect 3234 10792 3240 10804
rect 2731 10764 3240 10792
rect 2731 10761 2743 10764
rect 2685 10755 2743 10761
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 2130 10684 2136 10736
rect 2188 10724 2194 10736
rect 2188 10696 2544 10724
rect 2188 10684 2194 10696
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 2041 10659 2099 10665
rect 2041 10656 2053 10659
rect 1912 10628 2053 10656
rect 1912 10616 1918 10628
rect 2041 10625 2053 10628
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10656 2283 10659
rect 2314 10656 2320 10668
rect 2271 10628 2320 10656
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 2516 10665 2544 10696
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10625 2559 10659
rect 2501 10619 2559 10625
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4890 10656 4896 10668
rect 4387 10628 4896 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 9858 10656 9864 10668
rect 9819 10628 9864 10656
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 4614 10588 4620 10600
rect 4575 10560 4620 10588
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 10042 10520 10048 10532
rect 10003 10492 10048 10520
rect 10042 10480 10048 10492
rect 10100 10480 10106 10532
rect 1104 10362 10856 10384
rect 1104 10310 2582 10362
rect 2634 10310 2646 10362
rect 2698 10310 2710 10362
rect 2762 10310 2774 10362
rect 2826 10310 2838 10362
rect 2890 10310 5845 10362
rect 5897 10310 5909 10362
rect 5961 10310 5973 10362
rect 6025 10310 6037 10362
rect 6089 10310 6101 10362
rect 6153 10310 9109 10362
rect 9161 10310 9173 10362
rect 9225 10310 9237 10362
rect 9289 10310 9301 10362
rect 9353 10310 9365 10362
rect 9417 10310 10856 10362
rect 1104 10288 10856 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2222 10248 2228 10260
rect 1995 10220 2228 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 2038 10044 2044 10056
rect 1443 10016 2044 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 2038 10004 2044 10016
rect 2096 10004 2102 10056
rect 3970 10044 3976 10056
rect 3931 10016 3976 10044
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4614 10044 4620 10056
rect 4203 10016 4620 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 1026 9936 1032 9988
rect 1084 9976 1090 9988
rect 2222 9976 2228 9988
rect 1084 9948 2228 9976
rect 1084 9936 1090 9948
rect 2222 9936 2228 9948
rect 2280 9936 2286 9988
rect 4065 9911 4123 9917
rect 4065 9877 4077 9911
rect 4111 9908 4123 9911
rect 9858 9908 9864 9920
rect 4111 9880 9864 9908
rect 4111 9877 4123 9880
rect 4065 9871 4123 9877
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 1104 9818 10856 9840
rect 1104 9766 4213 9818
rect 4265 9766 4277 9818
rect 4329 9766 4341 9818
rect 4393 9766 4405 9818
rect 4457 9766 4469 9818
rect 4521 9766 7477 9818
rect 7529 9766 7541 9818
rect 7593 9766 7605 9818
rect 7657 9766 7669 9818
rect 7721 9766 7733 9818
rect 7785 9766 10856 9818
rect 1104 9744 10856 9766
rect 9858 9664 9864 9716
rect 9916 9664 9922 9716
rect 3694 9528 3700 9580
rect 3752 9568 3758 9580
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3752 9540 3985 9568
rect 3752 9528 3758 9540
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4614 9568 4620 9580
rect 4203 9540 4620 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 4890 9568 4896 9580
rect 4847 9540 4896 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 4890 9528 4896 9540
rect 4948 9528 4954 9580
rect 9876 9577 9904 9664
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 5074 9500 5080 9512
rect 5035 9472 5080 9500
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 10042 9432 10048 9444
rect 10003 9404 10048 9432
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 9858 9364 9864 9376
rect 4203 9336 9864 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 1104 9274 10856 9296
rect 1104 9222 2582 9274
rect 2634 9222 2646 9274
rect 2698 9222 2710 9274
rect 2762 9222 2774 9274
rect 2826 9222 2838 9274
rect 2890 9222 5845 9274
rect 5897 9222 5909 9274
rect 5961 9222 5973 9274
rect 6025 9222 6037 9274
rect 6089 9222 6101 9274
rect 6153 9222 9109 9274
rect 9161 9222 9173 9274
rect 9225 9222 9237 9274
rect 9289 9222 9301 9274
rect 9353 9222 9365 9274
rect 9417 9222 10856 9274
rect 1104 9200 10856 9222
rect 1104 8730 10856 8752
rect 1104 8678 4213 8730
rect 4265 8678 4277 8730
rect 4329 8678 4341 8730
rect 4393 8678 4405 8730
rect 4457 8678 4469 8730
rect 4521 8678 7477 8730
rect 7529 8678 7541 8730
rect 7593 8678 7605 8730
rect 7657 8678 7669 8730
rect 7721 8678 7733 8730
rect 7785 8678 10856 8730
rect 1104 8656 10856 8678
rect 9858 8480 9864 8492
rect 9819 8452 9864 8480
rect 9858 8440 9864 8452
rect 9916 8440 9922 8492
rect 10042 8344 10048 8356
rect 10003 8316 10048 8344
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 1104 8186 10856 8208
rect 1104 8134 2582 8186
rect 2634 8134 2646 8186
rect 2698 8134 2710 8186
rect 2762 8134 2774 8186
rect 2826 8134 2838 8186
rect 2890 8134 5845 8186
rect 5897 8134 5909 8186
rect 5961 8134 5973 8186
rect 6025 8134 6037 8186
rect 6089 8134 6101 8186
rect 6153 8134 9109 8186
rect 9161 8134 9173 8186
rect 9225 8134 9237 8186
rect 9289 8134 9301 8186
rect 9353 8134 9365 8186
rect 9417 8134 10856 8186
rect 1104 8112 10856 8134
rect 3878 7868 3884 7880
rect 3839 7840 3884 7868
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 4614 7868 4620 7880
rect 4111 7840 4620 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 3973 7735 4031 7741
rect 3973 7701 3985 7735
rect 4019 7732 4031 7735
rect 9858 7732 9864 7744
rect 4019 7704 9864 7732
rect 4019 7701 4031 7704
rect 3973 7695 4031 7701
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 1104 7642 10856 7664
rect 1104 7590 4213 7642
rect 4265 7590 4277 7642
rect 4329 7590 4341 7642
rect 4393 7590 4405 7642
rect 4457 7590 4469 7642
rect 4521 7590 7477 7642
rect 7529 7590 7541 7642
rect 7593 7590 7605 7642
rect 7657 7590 7669 7642
rect 7721 7590 7733 7642
rect 7785 7590 10856 7642
rect 1104 7568 10856 7590
rect 9858 7392 9864 7404
rect 9819 7364 9864 7392
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 10042 7256 10048 7268
rect 10003 7228 10048 7256
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 1104 7098 10856 7120
rect 1104 7046 2582 7098
rect 2634 7046 2646 7098
rect 2698 7046 2710 7098
rect 2762 7046 2774 7098
rect 2826 7046 2838 7098
rect 2890 7046 5845 7098
rect 5897 7046 5909 7098
rect 5961 7046 5973 7098
rect 6025 7046 6037 7098
rect 6089 7046 6101 7098
rect 6153 7046 9109 7098
rect 9161 7046 9173 7098
rect 9225 7046 9237 7098
rect 9289 7046 9301 7098
rect 9353 7046 9365 7098
rect 9417 7046 10856 7098
rect 1104 7024 10856 7046
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 3016 6752 4629 6780
rect 3016 6740 3022 6752
rect 4617 6749 4629 6752
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6780 4859 6783
rect 5074 6780 5080 6792
rect 4847 6752 5080 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 4709 6647 4767 6653
rect 4709 6613 4721 6647
rect 4755 6644 4767 6647
rect 9858 6644 9864 6656
rect 4755 6616 9864 6644
rect 4755 6613 4767 6616
rect 4709 6607 4767 6613
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 1104 6554 10856 6576
rect 1104 6502 4213 6554
rect 4265 6502 4277 6554
rect 4329 6502 4341 6554
rect 4393 6502 4405 6554
rect 4457 6502 4469 6554
rect 4521 6502 7477 6554
rect 7529 6502 7541 6554
rect 7593 6502 7605 6554
rect 7657 6502 7669 6554
rect 7721 6502 7733 6554
rect 7785 6502 10856 6554
rect 1104 6480 10856 6502
rect 2869 6443 2927 6449
rect 2869 6409 2881 6443
rect 2915 6440 2927 6443
rect 3878 6440 3884 6452
rect 2915 6412 3884 6440
rect 2915 6409 2927 6412
rect 2869 6403 2927 6409
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 2222 6372 2228 6384
rect 2135 6344 2228 6372
rect 2222 6332 2228 6344
rect 2280 6372 2286 6384
rect 2280 6344 4660 6372
rect 2280 6332 2286 6344
rect 1670 6264 1676 6316
rect 1728 6304 1734 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1728 6276 2145 6304
rect 1728 6264 1734 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 3142 6304 3148 6316
rect 2823 6276 3148 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 4632 6313 4660 6344
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 5074 6304 5080 6316
rect 4847 6276 5080 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 9858 6304 9864 6316
rect 9819 6276 9864 6304
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 3878 6128 3884 6180
rect 3936 6168 3942 6180
rect 6822 6168 6828 6180
rect 3936 6140 6828 6168
rect 3936 6128 3942 6140
rect 6822 6128 6828 6140
rect 6880 6128 6886 6180
rect 4801 6103 4859 6109
rect 4801 6069 4813 6103
rect 4847 6100 4859 6103
rect 9766 6100 9772 6112
rect 4847 6072 9772 6100
rect 4847 6069 4859 6072
rect 4801 6063 4859 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10042 6100 10048 6112
rect 10003 6072 10048 6100
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 1104 6010 10856 6032
rect 1104 5958 2582 6010
rect 2634 5958 2646 6010
rect 2698 5958 2710 6010
rect 2762 5958 2774 6010
rect 2826 5958 2838 6010
rect 2890 5958 5845 6010
rect 5897 5958 5909 6010
rect 5961 5958 5973 6010
rect 6025 5958 6037 6010
rect 6089 5958 6101 6010
rect 6153 5958 9109 6010
rect 9161 5958 9173 6010
rect 9225 5958 9237 6010
rect 9289 5958 9301 6010
rect 9353 5958 9365 6010
rect 9417 5958 10856 6010
rect 1104 5936 10856 5958
rect 1210 5856 1216 5908
rect 1268 5896 1274 5908
rect 2225 5899 2283 5905
rect 2225 5896 2237 5899
rect 1268 5868 2237 5896
rect 1268 5856 1274 5868
rect 1504 5760 1532 5868
rect 2225 5865 2237 5868
rect 2271 5865 2283 5899
rect 3878 5896 3884 5908
rect 2225 5859 2283 5865
rect 2332 5868 3884 5896
rect 1581 5831 1639 5837
rect 1581 5797 1593 5831
rect 1627 5828 1639 5831
rect 2332 5828 2360 5868
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 3973 5899 4031 5905
rect 3973 5865 3985 5899
rect 4019 5896 4031 5899
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 4019 5868 11069 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 1627 5800 2360 5828
rect 2869 5831 2927 5837
rect 1627 5797 1639 5800
rect 1581 5791 1639 5797
rect 2869 5797 2881 5831
rect 2915 5828 2927 5831
rect 3605 5831 3663 5837
rect 3605 5828 3617 5831
rect 2915 5800 3617 5828
rect 2915 5797 2927 5800
rect 2869 5791 2927 5797
rect 3605 5797 3617 5800
rect 3651 5828 3663 5831
rect 3651 5800 5304 5828
rect 3651 5797 3663 5800
rect 3605 5791 3663 5797
rect 1504 5732 4660 5760
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 1486 5692 1492 5704
rect 1443 5664 1492 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 1486 5652 1492 5664
rect 1544 5652 1550 5704
rect 2130 5692 2136 5704
rect 2091 5664 2136 5692
rect 2130 5652 2136 5664
rect 2188 5652 2194 5704
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 3050 5692 3056 5704
rect 2823 5664 3056 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 4632 5701 4660 5732
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 5074 5692 5080 5704
rect 4847 5664 5080 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 1504 5624 1532 5652
rect 3804 5624 3832 5655
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5276 5701 5304 5800
rect 5249 5695 5307 5701
rect 5249 5661 5261 5695
rect 5295 5661 5307 5695
rect 5249 5655 5307 5661
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 5408 5664 5457 5692
rect 5408 5652 5414 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 1504 5596 3832 5624
rect 4709 5627 4767 5633
rect 4709 5593 4721 5627
rect 4755 5624 4767 5627
rect 10965 5627 11023 5633
rect 10965 5624 10977 5627
rect 4755 5596 10977 5624
rect 4755 5593 4767 5596
rect 4709 5587 4767 5593
rect 10965 5593 10977 5596
rect 11011 5593 11023 5627
rect 10965 5587 11023 5593
rect 1118 5516 1124 5568
rect 1176 5556 1182 5568
rect 3605 5559 3663 5565
rect 3605 5556 3617 5559
rect 1176 5528 3617 5556
rect 1176 5516 1182 5528
rect 3605 5525 3617 5528
rect 3651 5525 3663 5559
rect 3605 5519 3663 5525
rect 5353 5559 5411 5565
rect 5353 5525 5365 5559
rect 5399 5556 5411 5559
rect 9858 5556 9864 5568
rect 5399 5528 9864 5556
rect 5399 5525 5411 5528
rect 5353 5519 5411 5525
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 1104 5466 10856 5488
rect 1104 5414 4213 5466
rect 4265 5414 4277 5466
rect 4329 5414 4341 5466
rect 4393 5414 4405 5466
rect 4457 5414 4469 5466
rect 4521 5414 7477 5466
rect 7529 5414 7541 5466
rect 7593 5414 7605 5466
rect 7657 5414 7669 5466
rect 7721 5414 7733 5466
rect 7785 5414 10856 5466
rect 1104 5392 10856 5414
rect 1302 5312 1308 5364
rect 1360 5352 1366 5364
rect 2225 5355 2283 5361
rect 2225 5352 2237 5355
rect 1360 5324 2237 5352
rect 1360 5312 1366 5324
rect 2225 5321 2237 5324
rect 2271 5321 2283 5355
rect 2225 5315 2283 5321
rect 2869 5355 2927 5361
rect 2869 5321 2881 5355
rect 2915 5352 2927 5355
rect 2958 5352 2964 5364
rect 2915 5324 2964 5352
rect 2915 5321 2927 5324
rect 2869 5315 2927 5321
rect 2240 5284 2268 5315
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 2240 5256 4660 5284
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 2133 5219 2191 5225
rect 2133 5216 2145 5219
rect 1636 5188 2145 5216
rect 1636 5176 1642 5188
rect 2133 5185 2145 5188
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5216 2835 5219
rect 2958 5216 2964 5228
rect 2823 5188 2964 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 4632 5225 4660 5256
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 5074 5216 5080 5228
rect 4847 5188 5080 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 9766 5176 9772 5228
rect 9824 5216 9830 5228
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9824 5188 9873 5216
rect 9824 5176 9830 5188
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 4798 5012 4804 5024
rect 4759 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 10042 5012 10048 5024
rect 10003 4984 10048 5012
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 1104 4922 10856 4944
rect 1104 4870 2582 4922
rect 2634 4870 2646 4922
rect 2698 4870 2710 4922
rect 2762 4870 2774 4922
rect 2826 4870 2838 4922
rect 2890 4870 5845 4922
rect 5897 4870 5909 4922
rect 5961 4870 5973 4922
rect 6025 4870 6037 4922
rect 6089 4870 6101 4922
rect 6153 4870 9109 4922
rect 9161 4870 9173 4922
rect 9225 4870 9237 4922
rect 9289 4870 9301 4922
rect 9353 4870 9365 4922
rect 9417 4870 10856 4922
rect 1104 4848 10856 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 3142 4808 3148 4820
rect 1627 4780 3148 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 1104 4378 10856 4400
rect 1104 4326 4213 4378
rect 4265 4326 4277 4378
rect 4329 4326 4341 4378
rect 4393 4326 4405 4378
rect 4457 4326 4469 4378
rect 4521 4326 7477 4378
rect 7529 4326 7541 4378
rect 7593 4326 7605 4378
rect 7657 4326 7669 4378
rect 7721 4326 7733 4378
rect 7785 4326 10856 4378
rect 1104 4304 10856 4326
rect 4798 4156 4804 4208
rect 4856 4196 4862 4208
rect 4856 4168 9904 4196
rect 4856 4156 4862 4168
rect 1210 4088 1216 4140
rect 1268 4128 1274 4140
rect 9876 4137 9904 4168
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 1268 4100 1409 4128
rect 1268 4088 1274 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 2958 3992 2964 4004
rect 1627 3964 2964 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 1104 3834 10856 3856
rect 1104 3782 2582 3834
rect 2634 3782 2646 3834
rect 2698 3782 2710 3834
rect 2762 3782 2774 3834
rect 2826 3782 2838 3834
rect 2890 3782 5845 3834
rect 5897 3782 5909 3834
rect 5961 3782 5973 3834
rect 6025 3782 6037 3834
rect 6089 3782 6101 3834
rect 6153 3782 9109 3834
rect 9161 3782 9173 3834
rect 9225 3782 9237 3834
rect 9289 3782 9301 3834
rect 9353 3782 9365 3834
rect 9417 3782 10856 3834
rect 1104 3760 10856 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 1670 3720 1676 3732
rect 1627 3692 1676 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 1670 3680 1676 3692
rect 1728 3680 1734 3732
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1360 3488 1409 3516
rect 1360 3476 1366 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 9858 3516 9864 3528
rect 9819 3488 9864 3516
rect 1397 3479 1455 3485
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 10042 3380 10048 3392
rect 10003 3352 10048 3380
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 1104 3290 10856 3312
rect 1104 3238 4213 3290
rect 4265 3238 4277 3290
rect 4329 3238 4341 3290
rect 4393 3238 4405 3290
rect 4457 3238 4469 3290
rect 4521 3238 7477 3290
rect 7529 3238 7541 3290
rect 7593 3238 7605 3290
rect 7657 3238 7669 3290
rect 7721 3238 7733 3290
rect 7785 3238 10856 3290
rect 1104 3216 10856 3238
rect 1578 3176 1584 3188
rect 1539 3148 1584 3176
rect 1578 3136 1584 3148
rect 1636 3136 1642 3188
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3040 9919 3043
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 9907 3012 10977 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 10045 2839 10103 2845
rect 10045 2805 10057 2839
rect 10091 2836 10103 2839
rect 10965 2839 11023 2845
rect 10965 2836 10977 2839
rect 10091 2808 10977 2836
rect 10091 2805 10103 2808
rect 10045 2799 10103 2805
rect 10965 2805 10977 2808
rect 11011 2805 11023 2839
rect 10965 2799 11023 2805
rect 1104 2746 10856 2768
rect 1104 2694 2582 2746
rect 2634 2694 2646 2746
rect 2698 2694 2710 2746
rect 2762 2694 2774 2746
rect 2826 2694 2838 2746
rect 2890 2694 5845 2746
rect 5897 2694 5909 2746
rect 5961 2694 5973 2746
rect 6025 2694 6037 2746
rect 6089 2694 6101 2746
rect 6153 2694 9109 2746
rect 9161 2694 9173 2746
rect 9225 2694 9237 2746
rect 9289 2694 9301 2746
rect 9353 2694 9365 2746
rect 9417 2694 10856 2746
rect 1104 2672 10856 2694
rect 1486 2592 1492 2644
rect 1544 2632 1550 2644
rect 1581 2635 1639 2641
rect 1581 2632 1593 2635
rect 1544 2604 1593 2632
rect 1544 2592 1550 2604
rect 1581 2601 1593 2604
rect 1627 2601 1639 2635
rect 1581 2595 1639 2601
rect 2130 2592 2136 2644
rect 2188 2632 2194 2644
rect 2225 2635 2283 2641
rect 2225 2632 2237 2635
rect 2188 2604 2237 2632
rect 2188 2592 2194 2604
rect 2225 2601 2237 2604
rect 2271 2601 2283 2635
rect 2225 2595 2283 2601
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 2958 2632 2964 2644
rect 2915 2604 2964 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 2038 2428 2044 2440
rect 1999 2400 2044 2428
rect 1397 2391 1455 2397
rect 2038 2388 2044 2400
rect 2096 2388 2102 2440
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 2774 2428 2780 2440
rect 2731 2400 2780 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2428 9919 2431
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 9907 2400 11069 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 10042 2292 10048 2304
rect 10003 2264 10048 2292
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 1104 2202 10856 2224
rect 1104 2150 4213 2202
rect 4265 2150 4277 2202
rect 4329 2150 4341 2202
rect 4393 2150 4405 2202
rect 4457 2150 4469 2202
rect 4521 2150 7477 2202
rect 7529 2150 7541 2202
rect 7593 2150 7605 2202
rect 7657 2150 7669 2202
rect 7721 2150 7733 2202
rect 7785 2150 10856 2202
rect 1104 2128 10856 2150
rect 10962 660 10968 672
rect 10923 632 10968 660
rect 10962 620 10968 632
rect 11020 620 11026 672
<< via1 >>
rect 10968 78251 11020 78260
rect 10968 78217 10977 78251
rect 10977 78217 11011 78251
rect 11011 78217 11020 78251
rect 10968 78208 11020 78217
rect 2582 77766 2634 77818
rect 2646 77766 2698 77818
rect 2710 77766 2762 77818
rect 2774 77766 2826 77818
rect 2838 77766 2890 77818
rect 5845 77766 5897 77818
rect 5909 77766 5961 77818
rect 5973 77766 6025 77818
rect 6037 77766 6089 77818
rect 6101 77766 6153 77818
rect 9109 77766 9161 77818
rect 9173 77766 9225 77818
rect 9237 77766 9289 77818
rect 9301 77766 9353 77818
rect 9365 77766 9417 77818
rect 1492 77460 1544 77512
rect 2044 77503 2096 77512
rect 2044 77469 2053 77503
rect 2053 77469 2087 77503
rect 2087 77469 2096 77503
rect 2044 77460 2096 77469
rect 2872 77503 2924 77512
rect 2872 77469 2881 77503
rect 2881 77469 2915 77503
rect 2915 77469 2924 77503
rect 2872 77460 2924 77469
rect 3976 77503 4028 77512
rect 3976 77469 3985 77503
rect 3985 77469 4019 77503
rect 4019 77469 4028 77503
rect 3976 77460 4028 77469
rect 9496 77503 9548 77512
rect 9496 77469 9505 77503
rect 9505 77469 9539 77503
rect 9539 77469 9548 77503
rect 9496 77460 9548 77469
rect 10140 77503 10192 77512
rect 10140 77469 10149 77503
rect 10149 77469 10183 77503
rect 10183 77469 10192 77503
rect 10140 77460 10192 77469
rect 1584 77367 1636 77376
rect 1584 77333 1593 77367
rect 1593 77333 1627 77367
rect 1627 77333 1636 77367
rect 1584 77324 1636 77333
rect 2136 77324 2188 77376
rect 2412 77324 2464 77376
rect 2872 77324 2924 77376
rect 5540 77324 5592 77376
rect 9680 77324 9732 77376
rect 4213 77222 4265 77274
rect 4277 77222 4329 77274
rect 4341 77222 4393 77274
rect 4405 77222 4457 77274
rect 4469 77222 4521 77274
rect 7477 77222 7529 77274
rect 7541 77222 7593 77274
rect 7605 77222 7657 77274
rect 7669 77222 7721 77274
rect 7733 77222 7785 77274
rect 1400 77027 1452 77036
rect 1400 76993 1409 77027
rect 1409 76993 1443 77027
rect 1443 76993 1452 77027
rect 1400 76984 1452 76993
rect 2044 77027 2096 77036
rect 2044 76993 2053 77027
rect 2053 76993 2087 77027
rect 2087 76993 2096 77027
rect 2044 76984 2096 76993
rect 2964 76984 3016 77036
rect 1676 76780 1728 76832
rect 2320 76780 2372 76832
rect 2504 76780 2556 76832
rect 9956 76823 10008 76832
rect 9956 76789 9965 76823
rect 9965 76789 9999 76823
rect 9999 76789 10008 76823
rect 9956 76780 10008 76789
rect 2582 76678 2634 76730
rect 2646 76678 2698 76730
rect 2710 76678 2762 76730
rect 2774 76678 2826 76730
rect 2838 76678 2890 76730
rect 5845 76678 5897 76730
rect 5909 76678 5961 76730
rect 5973 76678 6025 76730
rect 6037 76678 6089 76730
rect 6101 76678 6153 76730
rect 9109 76678 9161 76730
rect 9173 76678 9225 76730
rect 9237 76678 9289 76730
rect 9301 76678 9353 76730
rect 9365 76678 9417 76730
rect 1308 76372 1360 76424
rect 3056 76440 3108 76492
rect 3148 76372 3200 76424
rect 10140 76415 10192 76424
rect 10140 76381 10149 76415
rect 10149 76381 10183 76415
rect 10183 76381 10192 76415
rect 10140 76372 10192 76381
rect 3516 76304 3568 76356
rect 2044 76279 2096 76288
rect 2044 76245 2053 76279
rect 2053 76245 2087 76279
rect 2087 76245 2096 76279
rect 2044 76236 2096 76245
rect 3148 76236 3200 76288
rect 9772 76236 9824 76288
rect 4213 76134 4265 76186
rect 4277 76134 4329 76186
rect 4341 76134 4393 76186
rect 4405 76134 4457 76186
rect 4469 76134 4521 76186
rect 7477 76134 7529 76186
rect 7541 76134 7593 76186
rect 7605 76134 7657 76186
rect 7669 76134 7721 76186
rect 7733 76134 7785 76186
rect 1860 76032 1912 76084
rect 1952 76032 2004 76084
rect 1400 75939 1452 75948
rect 1400 75905 1409 75939
rect 1409 75905 1443 75939
rect 1443 75905 1452 75939
rect 1400 75896 1452 75905
rect 1492 75896 1544 75948
rect 1676 75896 1728 75948
rect 2228 75939 2280 75948
rect 2228 75905 2237 75939
rect 2237 75905 2271 75939
rect 2271 75905 2280 75939
rect 2228 75896 2280 75905
rect 2582 75590 2634 75642
rect 2646 75590 2698 75642
rect 2710 75590 2762 75642
rect 2774 75590 2826 75642
rect 2838 75590 2890 75642
rect 5845 75590 5897 75642
rect 5909 75590 5961 75642
rect 5973 75590 6025 75642
rect 6037 75590 6089 75642
rect 6101 75590 6153 75642
rect 9109 75590 9161 75642
rect 9173 75590 9225 75642
rect 9237 75590 9289 75642
rect 9301 75590 9353 75642
rect 9365 75590 9417 75642
rect 1124 75420 1176 75472
rect 940 75216 992 75268
rect 2044 75327 2096 75336
rect 2044 75293 2053 75327
rect 2053 75293 2087 75327
rect 2087 75293 2096 75327
rect 2320 75327 2372 75336
rect 2044 75284 2096 75293
rect 2320 75293 2329 75327
rect 2329 75293 2363 75327
rect 2363 75293 2372 75327
rect 2320 75284 2372 75293
rect 2780 75327 2832 75336
rect 2780 75293 2789 75327
rect 2789 75293 2823 75327
rect 2823 75293 2832 75327
rect 2780 75284 2832 75293
rect 9956 75284 10008 75336
rect 10140 75327 10192 75336
rect 10140 75293 10149 75327
rect 10149 75293 10183 75327
rect 10183 75293 10192 75327
rect 10140 75284 10192 75293
rect 2596 75148 2648 75200
rect 4620 75148 4672 75200
rect 9864 75148 9916 75200
rect 4213 75046 4265 75098
rect 4277 75046 4329 75098
rect 4341 75046 4393 75098
rect 4405 75046 4457 75098
rect 4469 75046 4521 75098
rect 7477 75046 7529 75098
rect 7541 75046 7593 75098
rect 7605 75046 7657 75098
rect 7669 75046 7721 75098
rect 7733 75046 7785 75098
rect 940 74808 992 74860
rect 9680 74944 9732 74996
rect 2872 74876 2924 74928
rect 3148 74919 3200 74928
rect 3148 74885 3157 74919
rect 3157 74885 3191 74919
rect 3191 74885 3200 74919
rect 3148 74876 3200 74885
rect 5540 74876 5592 74928
rect 2320 74851 2372 74860
rect 2320 74817 2329 74851
rect 2329 74817 2363 74851
rect 2363 74817 2372 74851
rect 2320 74808 2372 74817
rect 2596 74808 2648 74860
rect 5172 74808 5224 74860
rect 3700 74672 3752 74724
rect 2964 74604 3016 74656
rect 2582 74502 2634 74554
rect 2646 74502 2698 74554
rect 2710 74502 2762 74554
rect 2774 74502 2826 74554
rect 2838 74502 2890 74554
rect 5845 74502 5897 74554
rect 5909 74502 5961 74554
rect 5973 74502 6025 74554
rect 6037 74502 6089 74554
rect 6101 74502 6153 74554
rect 9109 74502 9161 74554
rect 9173 74502 9225 74554
rect 9237 74502 9289 74554
rect 9301 74502 9353 74554
rect 9365 74502 9417 74554
rect 8300 74332 8352 74384
rect 2596 74264 2648 74316
rect 3516 74264 3568 74316
rect 1308 74196 1360 74248
rect 2320 74239 2372 74248
rect 2320 74205 2369 74239
rect 2369 74205 2372 74239
rect 2320 74196 2372 74205
rect 2504 74239 2556 74248
rect 2504 74205 2513 74239
rect 2513 74205 2547 74239
rect 2547 74205 2556 74239
rect 2780 74239 2832 74248
rect 2504 74196 2556 74205
rect 2780 74205 2789 74239
rect 2789 74205 2823 74239
rect 2823 74205 2832 74239
rect 2780 74196 2832 74205
rect 2872 74196 2924 74248
rect 10140 74239 10192 74248
rect 10140 74205 10149 74239
rect 10149 74205 10183 74239
rect 10183 74205 10192 74239
rect 10140 74196 10192 74205
rect 9772 74128 9824 74180
rect 1676 74060 1728 74112
rect 3976 74060 4028 74112
rect 9956 74103 10008 74112
rect 9956 74069 9965 74103
rect 9965 74069 9999 74103
rect 9999 74069 10008 74103
rect 9956 74060 10008 74069
rect 4213 73958 4265 74010
rect 4277 73958 4329 74010
rect 4341 73958 4393 74010
rect 4405 73958 4457 74010
rect 4469 73958 4521 74010
rect 7477 73958 7529 74010
rect 7541 73958 7593 74010
rect 7605 73958 7657 74010
rect 7669 73958 7721 74010
rect 7733 73958 7785 74010
rect 2412 73856 2464 73908
rect 9864 73788 9916 73840
rect 1400 73763 1452 73772
rect 1400 73729 1409 73763
rect 1409 73729 1443 73763
rect 1443 73729 1452 73763
rect 1400 73720 1452 73729
rect 2320 73763 2372 73772
rect 2320 73729 2369 73763
rect 2369 73729 2372 73763
rect 2780 73763 2832 73772
rect 2320 73720 2372 73729
rect 2780 73729 2789 73763
rect 2789 73729 2823 73763
rect 2823 73729 2832 73763
rect 2780 73720 2832 73729
rect 3056 73720 3108 73772
rect 2412 73584 2464 73636
rect 4988 73516 5040 73568
rect 2582 73414 2634 73466
rect 2646 73414 2698 73466
rect 2710 73414 2762 73466
rect 2774 73414 2826 73466
rect 2838 73414 2890 73466
rect 5845 73414 5897 73466
rect 5909 73414 5961 73466
rect 5973 73414 6025 73466
rect 6037 73414 6089 73466
rect 6101 73414 6153 73466
rect 9109 73414 9161 73466
rect 9173 73414 9225 73466
rect 9237 73414 9289 73466
rect 9301 73414 9353 73466
rect 9365 73414 9417 73466
rect 1308 73108 1360 73160
rect 2320 73151 2372 73160
rect 2320 73117 2369 73151
rect 2369 73117 2372 73151
rect 2320 73108 2372 73117
rect 3056 73108 3108 73160
rect 5540 73108 5592 73160
rect 2136 73040 2188 73092
rect 9956 73108 10008 73160
rect 10140 73151 10192 73160
rect 10140 73117 10149 73151
rect 10149 73117 10183 73151
rect 10183 73117 10192 73151
rect 10140 73108 10192 73117
rect 3148 72972 3200 73024
rect 8392 72972 8444 73024
rect 4213 72870 4265 72922
rect 4277 72870 4329 72922
rect 4341 72870 4393 72922
rect 4405 72870 4457 72922
rect 4469 72870 4521 72922
rect 7477 72870 7529 72922
rect 7541 72870 7593 72922
rect 7605 72870 7657 72922
rect 7669 72870 7721 72922
rect 7733 72870 7785 72922
rect 1860 72768 1912 72820
rect 2136 72768 2188 72820
rect 1216 72632 1268 72684
rect 2044 72675 2096 72684
rect 2044 72641 2053 72675
rect 2053 72641 2087 72675
rect 2087 72641 2096 72675
rect 2044 72632 2096 72641
rect 1768 72428 1820 72480
rect 1860 72428 1912 72480
rect 2582 72326 2634 72378
rect 2646 72326 2698 72378
rect 2710 72326 2762 72378
rect 2774 72326 2826 72378
rect 2838 72326 2890 72378
rect 5845 72326 5897 72378
rect 5909 72326 5961 72378
rect 5973 72326 6025 72378
rect 6037 72326 6089 72378
rect 6101 72326 6153 72378
rect 9109 72326 9161 72378
rect 9173 72326 9225 72378
rect 9237 72326 9289 72378
rect 9301 72326 9353 72378
rect 9365 72326 9417 72378
rect 1032 72156 1084 72208
rect 1400 72063 1452 72072
rect 1400 72029 1409 72063
rect 1409 72029 1443 72063
rect 1443 72029 1452 72063
rect 1400 72020 1452 72029
rect 1492 72020 1544 72072
rect 2044 72020 2096 72072
rect 2320 72063 2372 72072
rect 2320 72029 2369 72063
rect 2369 72029 2372 72063
rect 2320 72020 2372 72029
rect 3056 72020 3108 72072
rect 10140 72063 10192 72072
rect 10140 72029 10149 72063
rect 10149 72029 10183 72063
rect 10183 72029 10192 72063
rect 10140 72020 10192 72029
rect 1492 71884 1544 71936
rect 2228 71952 2280 72004
rect 8392 71952 8444 72004
rect 2320 71884 2372 71936
rect 9956 71927 10008 71936
rect 9956 71893 9965 71927
rect 9965 71893 9999 71927
rect 9999 71893 10008 71927
rect 9956 71884 10008 71893
rect 4213 71782 4265 71834
rect 4277 71782 4329 71834
rect 4341 71782 4393 71834
rect 4405 71782 4457 71834
rect 4469 71782 4521 71834
rect 7477 71782 7529 71834
rect 7541 71782 7593 71834
rect 7605 71782 7657 71834
rect 7669 71782 7721 71834
rect 7733 71782 7785 71834
rect 1584 71612 1636 71664
rect 9956 71612 10008 71664
rect 1308 71544 1360 71596
rect 2044 71544 2096 71596
rect 3056 71544 3108 71596
rect 1584 71383 1636 71392
rect 1584 71349 1593 71383
rect 1593 71349 1627 71383
rect 1627 71349 1636 71383
rect 1584 71340 1636 71349
rect 3240 71340 3292 71392
rect 2582 71238 2634 71290
rect 2646 71238 2698 71290
rect 2710 71238 2762 71290
rect 2774 71238 2826 71290
rect 2838 71238 2890 71290
rect 5845 71238 5897 71290
rect 5909 71238 5961 71290
rect 5973 71238 6025 71290
rect 6037 71238 6089 71290
rect 6101 71238 6153 71290
rect 9109 71238 9161 71290
rect 9173 71238 9225 71290
rect 9237 71238 9289 71290
rect 9301 71238 9353 71290
rect 9365 71238 9417 71290
rect 388 71068 440 71120
rect 2320 71068 2372 71120
rect 2596 71068 2648 71120
rect 1400 70975 1452 70984
rect 1400 70941 1409 70975
rect 1409 70941 1443 70975
rect 1443 70941 1452 70975
rect 1400 70932 1452 70941
rect 2320 70932 2372 70984
rect 2780 70932 2832 70984
rect 10140 70975 10192 70984
rect 10140 70941 10149 70975
rect 10149 70941 10183 70975
rect 10183 70941 10192 70975
rect 10140 70932 10192 70941
rect 1952 70864 2004 70916
rect 9864 70864 9916 70916
rect 2228 70796 2280 70848
rect 9956 70839 10008 70848
rect 9956 70805 9965 70839
rect 9965 70805 9999 70839
rect 9999 70805 10008 70839
rect 9956 70796 10008 70805
rect 4213 70694 4265 70746
rect 4277 70694 4329 70746
rect 4341 70694 4393 70746
rect 4405 70694 4457 70746
rect 4469 70694 4521 70746
rect 7477 70694 7529 70746
rect 7541 70694 7593 70746
rect 7605 70694 7657 70746
rect 7669 70694 7721 70746
rect 7733 70694 7785 70746
rect 1400 70524 1452 70576
rect 2596 70524 2648 70576
rect 9956 70524 10008 70576
rect 1216 70388 1268 70440
rect 1952 70388 2004 70440
rect 2320 70388 2372 70440
rect 3332 70456 3384 70508
rect 5264 70388 5316 70440
rect 2582 70150 2634 70202
rect 2646 70150 2698 70202
rect 2710 70150 2762 70202
rect 2774 70150 2826 70202
rect 2838 70150 2890 70202
rect 5845 70150 5897 70202
rect 5909 70150 5961 70202
rect 5973 70150 6025 70202
rect 6037 70150 6089 70202
rect 6101 70150 6153 70202
rect 9109 70150 9161 70202
rect 9173 70150 9225 70202
rect 9237 70150 9289 70202
rect 9301 70150 9353 70202
rect 9365 70150 9417 70202
rect 9864 70048 9916 70100
rect 1400 69980 1452 70032
rect 1584 69980 1636 70032
rect 848 69912 900 69964
rect 1400 69887 1452 69896
rect 1400 69853 1409 69887
rect 1409 69853 1443 69887
rect 1443 69853 1452 69887
rect 1400 69844 1452 69853
rect 2872 69887 2924 69896
rect 2872 69853 2881 69887
rect 2881 69853 2915 69887
rect 2915 69853 2924 69887
rect 2872 69844 2924 69853
rect 10140 69887 10192 69896
rect 10140 69853 10149 69887
rect 10149 69853 10183 69887
rect 10183 69853 10192 69887
rect 10140 69844 10192 69853
rect 2228 69708 2280 69760
rect 4213 69606 4265 69658
rect 4277 69606 4329 69658
rect 4341 69606 4393 69658
rect 4405 69606 4457 69658
rect 4469 69606 4521 69658
rect 7477 69606 7529 69658
rect 7541 69606 7593 69658
rect 7605 69606 7657 69658
rect 7669 69606 7721 69658
rect 7733 69606 7785 69658
rect 2044 69436 2096 69488
rect 3056 69436 3108 69488
rect 1308 69300 1360 69352
rect 2044 69300 2096 69352
rect 3056 69300 3108 69352
rect 3424 69300 3476 69352
rect 2582 69062 2634 69114
rect 2646 69062 2698 69114
rect 2710 69062 2762 69114
rect 2774 69062 2826 69114
rect 2838 69062 2890 69114
rect 5845 69062 5897 69114
rect 5909 69062 5961 69114
rect 5973 69062 6025 69114
rect 6037 69062 6089 69114
rect 6101 69062 6153 69114
rect 9109 69062 9161 69114
rect 9173 69062 9225 69114
rect 9237 69062 9289 69114
rect 9301 69062 9353 69114
rect 9365 69062 9417 69114
rect 1584 68892 1636 68944
rect 2320 68892 2372 68944
rect 3884 68935 3936 68944
rect 3884 68901 3893 68935
rect 3893 68901 3927 68935
rect 3927 68901 3936 68935
rect 3884 68892 3936 68901
rect 1400 68799 1452 68808
rect 1400 68765 1409 68799
rect 1409 68765 1443 68799
rect 1443 68765 1452 68799
rect 1400 68756 1452 68765
rect 1584 68756 1636 68808
rect 3332 68756 3384 68808
rect 4712 68756 4764 68808
rect 10140 68799 10192 68808
rect 10140 68765 10149 68799
rect 10149 68765 10183 68799
rect 10183 68765 10192 68799
rect 10140 68756 10192 68765
rect 2504 68688 2556 68740
rect 1768 68620 1820 68672
rect 2596 68620 2648 68672
rect 4213 68518 4265 68570
rect 4277 68518 4329 68570
rect 4341 68518 4393 68570
rect 4405 68518 4457 68570
rect 4469 68518 4521 68570
rect 7477 68518 7529 68570
rect 7541 68518 7593 68570
rect 7605 68518 7657 68570
rect 7669 68518 7721 68570
rect 7733 68518 7785 68570
rect 1860 68416 1912 68468
rect 2228 68416 2280 68468
rect 1492 68212 1544 68264
rect 1492 68119 1544 68128
rect 1492 68085 1501 68119
rect 1501 68085 1535 68119
rect 1535 68085 1544 68119
rect 1492 68076 1544 68085
rect 1768 68076 1820 68128
rect 2320 68280 2372 68332
rect 3056 68348 3108 68400
rect 3516 68348 3568 68400
rect 4620 68348 4672 68400
rect 3332 68280 3384 68332
rect 4344 68323 4396 68332
rect 4344 68289 4353 68323
rect 4353 68289 4387 68323
rect 4387 68289 4396 68323
rect 4344 68280 4396 68289
rect 4712 68280 4764 68332
rect 9956 68144 10008 68196
rect 2136 68076 2188 68128
rect 8392 68076 8444 68128
rect 2582 67974 2634 68026
rect 2646 67974 2698 68026
rect 2710 67974 2762 68026
rect 2774 67974 2826 68026
rect 2838 67974 2890 68026
rect 5845 67974 5897 68026
rect 5909 67974 5961 68026
rect 5973 67974 6025 68026
rect 6037 67974 6089 68026
rect 6101 67974 6153 68026
rect 9109 67974 9161 68026
rect 9173 67974 9225 68026
rect 9237 67974 9289 68026
rect 9301 67974 9353 68026
rect 9365 67974 9417 68026
rect 1492 67872 1544 67924
rect 4344 67872 4396 67924
rect 6920 67804 6972 67856
rect 2320 67736 2372 67788
rect 3424 67736 3476 67788
rect 3608 67736 3660 67788
rect 1676 67643 1728 67652
rect 1676 67609 1685 67643
rect 1685 67609 1719 67643
rect 1719 67609 1728 67643
rect 1676 67600 1728 67609
rect 4712 67600 4764 67652
rect 10140 67532 10192 67584
rect 4213 67430 4265 67482
rect 4277 67430 4329 67482
rect 4341 67430 4393 67482
rect 4405 67430 4457 67482
rect 4469 67430 4521 67482
rect 7477 67430 7529 67482
rect 7541 67430 7593 67482
rect 7605 67430 7657 67482
rect 7669 67430 7721 67482
rect 7733 67430 7785 67482
rect 1400 67235 1452 67244
rect 1400 67201 1409 67235
rect 1409 67201 1443 67235
rect 1443 67201 1452 67235
rect 1400 67192 1452 67201
rect 1676 66988 1728 67040
rect 2582 66886 2634 66938
rect 2646 66886 2698 66938
rect 2710 66886 2762 66938
rect 2774 66886 2826 66938
rect 2838 66886 2890 66938
rect 5845 66886 5897 66938
rect 5909 66886 5961 66938
rect 5973 66886 6025 66938
rect 6037 66886 6089 66938
rect 6101 66886 6153 66938
rect 9109 66886 9161 66938
rect 9173 66886 9225 66938
rect 9237 66886 9289 66938
rect 9301 66886 9353 66938
rect 9365 66886 9417 66938
rect 1400 66512 1452 66564
rect 2780 66512 2832 66564
rect 664 66444 716 66496
rect 3424 66444 3476 66496
rect 4213 66342 4265 66394
rect 4277 66342 4329 66394
rect 4341 66342 4393 66394
rect 4405 66342 4457 66394
rect 4469 66342 4521 66394
rect 7477 66342 7529 66394
rect 7541 66342 7593 66394
rect 7605 66342 7657 66394
rect 7669 66342 7721 66394
rect 7733 66342 7785 66394
rect 1952 66240 2004 66292
rect 2136 66240 2188 66292
rect 9956 66283 10008 66292
rect 9956 66249 9965 66283
rect 9965 66249 9999 66283
rect 9999 66249 10008 66283
rect 9956 66240 10008 66249
rect 1952 66147 2004 66156
rect 1952 66113 1961 66147
rect 1961 66113 1995 66147
rect 1995 66113 2004 66147
rect 1952 66104 2004 66113
rect 4068 66104 4120 66156
rect 10140 66147 10192 66156
rect 10140 66113 10149 66147
rect 10149 66113 10183 66147
rect 10183 66113 10192 66147
rect 10140 66104 10192 66113
rect 8484 65968 8536 66020
rect 3148 65900 3200 65952
rect 2582 65798 2634 65850
rect 2646 65798 2698 65850
rect 2710 65798 2762 65850
rect 2774 65798 2826 65850
rect 2838 65798 2890 65850
rect 5845 65798 5897 65850
rect 5909 65798 5961 65850
rect 5973 65798 6025 65850
rect 6037 65798 6089 65850
rect 6101 65798 6153 65850
rect 9109 65798 9161 65850
rect 9173 65798 9225 65850
rect 9237 65798 9289 65850
rect 9301 65798 9353 65850
rect 9365 65798 9417 65850
rect 2320 65628 2372 65680
rect 3056 65628 3108 65680
rect 3792 65492 3844 65544
rect 756 65424 808 65476
rect 1952 65467 2004 65476
rect 1952 65433 1961 65467
rect 1961 65433 1995 65467
rect 1995 65433 2004 65467
rect 1952 65424 2004 65433
rect 3056 65356 3108 65408
rect 4213 65254 4265 65306
rect 4277 65254 4329 65306
rect 4341 65254 4393 65306
rect 4405 65254 4457 65306
rect 4469 65254 4521 65306
rect 7477 65254 7529 65306
rect 7541 65254 7593 65306
rect 7605 65254 7657 65306
rect 7669 65254 7721 65306
rect 7733 65254 7785 65306
rect 5080 65084 5132 65136
rect 1952 65016 2004 65068
rect 2320 65016 2372 65068
rect 3516 65016 3568 65068
rect 10140 65059 10192 65068
rect 10140 65025 10149 65059
rect 10149 65025 10183 65059
rect 10183 65025 10192 65059
rect 10140 65016 10192 65025
rect 1492 64923 1544 64932
rect 1492 64889 1501 64923
rect 1501 64889 1535 64923
rect 1535 64889 1544 64923
rect 1492 64880 1544 64889
rect 940 64812 992 64864
rect 2320 64812 2372 64864
rect 9956 64855 10008 64864
rect 9956 64821 9965 64855
rect 9965 64821 9999 64855
rect 9999 64821 10008 64855
rect 9956 64812 10008 64821
rect 2582 64710 2634 64762
rect 2646 64710 2698 64762
rect 2710 64710 2762 64762
rect 2774 64710 2826 64762
rect 2838 64710 2890 64762
rect 5845 64710 5897 64762
rect 5909 64710 5961 64762
rect 5973 64710 6025 64762
rect 6037 64710 6089 64762
rect 6101 64710 6153 64762
rect 9109 64710 9161 64762
rect 9173 64710 9225 64762
rect 9237 64710 9289 64762
rect 9301 64710 9353 64762
rect 9365 64710 9417 64762
rect 20 64540 72 64592
rect 2320 64447 2372 64456
rect 2320 64413 2324 64447
rect 2324 64413 2358 64447
rect 2358 64413 2372 64447
rect 2320 64404 2372 64413
rect 3976 64472 4028 64524
rect 2780 64404 2832 64456
rect 3332 64404 3384 64456
rect 9956 64336 10008 64388
rect 3976 64311 4028 64320
rect 3976 64277 3985 64311
rect 3985 64277 4019 64311
rect 4019 64277 4028 64311
rect 3976 64268 4028 64277
rect 4213 64166 4265 64218
rect 4277 64166 4329 64218
rect 4341 64166 4393 64218
rect 4405 64166 4457 64218
rect 4469 64166 4521 64218
rect 7477 64166 7529 64218
rect 7541 64166 7593 64218
rect 7605 64166 7657 64218
rect 7669 64166 7721 64218
rect 7733 64166 7785 64218
rect 1400 63996 1452 64048
rect 940 63928 992 63980
rect 2320 63971 2372 63980
rect 2320 63937 2369 63971
rect 2369 63937 2372 63971
rect 2320 63928 2372 63937
rect 2780 63971 2832 63980
rect 2780 63937 2789 63971
rect 2789 63937 2823 63971
rect 2823 63937 2832 63971
rect 2780 63928 2832 63937
rect 3056 63928 3108 63980
rect 10140 63971 10192 63980
rect 10140 63937 10149 63971
rect 10149 63937 10183 63971
rect 10183 63937 10192 63971
rect 10140 63928 10192 63937
rect 1400 63724 1452 63776
rect 6736 63724 6788 63776
rect 2582 63622 2634 63674
rect 2646 63622 2698 63674
rect 2710 63622 2762 63674
rect 2774 63622 2826 63674
rect 2838 63622 2890 63674
rect 5845 63622 5897 63674
rect 5909 63622 5961 63674
rect 5973 63622 6025 63674
rect 6037 63622 6089 63674
rect 6101 63622 6153 63674
rect 9109 63622 9161 63674
rect 9173 63622 9225 63674
rect 9237 63622 9289 63674
rect 9301 63622 9353 63674
rect 9365 63622 9417 63674
rect 3516 63384 3568 63436
rect 5724 63316 5776 63368
rect 7380 63248 7432 63300
rect 1492 63223 1544 63232
rect 1492 63189 1501 63223
rect 1501 63189 1535 63223
rect 1535 63189 1544 63223
rect 1492 63180 1544 63189
rect 2320 63180 2372 63232
rect 3976 63223 4028 63232
rect 3976 63189 3985 63223
rect 3985 63189 4019 63223
rect 4019 63189 4028 63223
rect 3976 63180 4028 63189
rect 4213 63078 4265 63130
rect 4277 63078 4329 63130
rect 4341 63078 4393 63130
rect 4405 63078 4457 63130
rect 4469 63078 4521 63130
rect 7477 63078 7529 63130
rect 7541 63078 7593 63130
rect 7605 63078 7657 63130
rect 7669 63078 7721 63130
rect 7733 63078 7785 63130
rect 2412 62976 2464 63028
rect 3056 62840 3108 62892
rect 10140 62883 10192 62892
rect 10140 62849 10149 62883
rect 10149 62849 10183 62883
rect 10183 62849 10192 62883
rect 10140 62840 10192 62849
rect 2320 62772 2372 62824
rect 3148 62772 3200 62824
rect 3608 62772 3660 62824
rect 8576 62636 8628 62688
rect 2582 62534 2634 62586
rect 2646 62534 2698 62586
rect 2710 62534 2762 62586
rect 2774 62534 2826 62586
rect 2838 62534 2890 62586
rect 5845 62534 5897 62586
rect 5909 62534 5961 62586
rect 5973 62534 6025 62586
rect 6037 62534 6089 62586
rect 6101 62534 6153 62586
rect 9109 62534 9161 62586
rect 9173 62534 9225 62586
rect 9237 62534 9289 62586
rect 9301 62534 9353 62586
rect 9365 62534 9417 62586
rect 4620 62364 4672 62416
rect 1400 62092 1452 62144
rect 2320 62271 2372 62280
rect 2320 62237 2369 62271
rect 2369 62237 2372 62271
rect 2320 62228 2372 62237
rect 3056 62228 3108 62280
rect 1952 62160 2004 62212
rect 9956 62160 10008 62212
rect 7288 62092 7340 62144
rect 4213 61990 4265 62042
rect 4277 61990 4329 62042
rect 4341 61990 4393 62042
rect 4405 61990 4457 62042
rect 4469 61990 4521 62042
rect 7477 61990 7529 62042
rect 7541 61990 7593 62042
rect 7605 61990 7657 62042
rect 7669 61990 7721 62042
rect 7733 61990 7785 62042
rect 2228 61820 2280 61872
rect 296 61752 348 61804
rect 2320 61795 2372 61804
rect 2320 61761 2369 61795
rect 2369 61761 2372 61795
rect 2320 61752 2372 61761
rect 3056 61752 3108 61804
rect 10140 61795 10192 61804
rect 10140 61761 10149 61795
rect 10149 61761 10183 61795
rect 10183 61761 10192 61795
rect 10140 61752 10192 61761
rect 1492 61591 1544 61600
rect 1492 61557 1501 61591
rect 1501 61557 1535 61591
rect 1535 61557 1544 61591
rect 1492 61548 1544 61557
rect 8668 61548 8720 61600
rect 2582 61446 2634 61498
rect 2646 61446 2698 61498
rect 2710 61446 2762 61498
rect 2774 61446 2826 61498
rect 2838 61446 2890 61498
rect 5845 61446 5897 61498
rect 5909 61446 5961 61498
rect 5973 61446 6025 61498
rect 6037 61446 6089 61498
rect 6101 61446 6153 61498
rect 9109 61446 9161 61498
rect 9173 61446 9225 61498
rect 9237 61446 9289 61498
rect 9301 61446 9353 61498
rect 9365 61446 9417 61498
rect 2228 61387 2280 61396
rect 2228 61353 2237 61387
rect 2237 61353 2271 61387
rect 2271 61353 2280 61387
rect 2228 61344 2280 61353
rect 4896 61140 4948 61192
rect 5632 61072 5684 61124
rect 1400 61004 1452 61056
rect 4213 60902 4265 60954
rect 4277 60902 4329 60954
rect 4341 60902 4393 60954
rect 4405 60902 4457 60954
rect 4469 60902 4521 60954
rect 7477 60902 7529 60954
rect 7541 60902 7593 60954
rect 7605 60902 7657 60954
rect 7669 60902 7721 60954
rect 7733 60902 7785 60954
rect 1676 60800 1728 60852
rect 9956 60843 10008 60852
rect 9956 60809 9965 60843
rect 9965 60809 9999 60843
rect 9999 60809 10008 60843
rect 9956 60800 10008 60809
rect 480 60664 532 60716
rect 10140 60707 10192 60716
rect 10140 60673 10149 60707
rect 10149 60673 10183 60707
rect 10183 60673 10192 60707
rect 10140 60664 10192 60673
rect 1492 60503 1544 60512
rect 1492 60469 1501 60503
rect 1501 60469 1535 60503
rect 1535 60469 1544 60503
rect 1492 60460 1544 60469
rect 2582 60358 2634 60410
rect 2646 60358 2698 60410
rect 2710 60358 2762 60410
rect 2774 60358 2826 60410
rect 2838 60358 2890 60410
rect 5845 60358 5897 60410
rect 5909 60358 5961 60410
rect 5973 60358 6025 60410
rect 6037 60358 6089 60410
rect 6101 60358 6153 60410
rect 9109 60358 9161 60410
rect 9173 60358 9225 60410
rect 9237 60358 9289 60410
rect 9301 60358 9353 60410
rect 9365 60358 9417 60410
rect 6276 60052 6328 60104
rect 1400 59916 1452 59968
rect 4213 59814 4265 59866
rect 4277 59814 4329 59866
rect 4341 59814 4393 59866
rect 4405 59814 4457 59866
rect 4469 59814 4521 59866
rect 7477 59814 7529 59866
rect 7541 59814 7593 59866
rect 7605 59814 7657 59866
rect 7669 59814 7721 59866
rect 7733 59814 7785 59866
rect 572 59576 624 59628
rect 5356 59576 5408 59628
rect 10140 59619 10192 59628
rect 10140 59585 10149 59619
rect 10149 59585 10183 59619
rect 10183 59585 10192 59619
rect 10140 59576 10192 59585
rect 2228 59483 2280 59492
rect 2228 59449 2237 59483
rect 2237 59449 2271 59483
rect 2271 59449 2280 59483
rect 2228 59440 2280 59449
rect 1492 59415 1544 59424
rect 1492 59381 1501 59415
rect 1501 59381 1535 59415
rect 1535 59381 1544 59415
rect 1492 59372 1544 59381
rect 9956 59415 10008 59424
rect 9956 59381 9965 59415
rect 9965 59381 9999 59415
rect 9999 59381 10008 59415
rect 9956 59372 10008 59381
rect 2582 59270 2634 59322
rect 2646 59270 2698 59322
rect 2710 59270 2762 59322
rect 2774 59270 2826 59322
rect 2838 59270 2890 59322
rect 5845 59270 5897 59322
rect 5909 59270 5961 59322
rect 5973 59270 6025 59322
rect 6037 59270 6089 59322
rect 6101 59270 6153 59322
rect 9109 59270 9161 59322
rect 9173 59270 9225 59322
rect 9237 59270 9289 59322
rect 9301 59270 9353 59322
rect 9365 59270 9417 59322
rect 3884 59100 3936 59152
rect 2320 59032 2372 59084
rect 2228 58964 2280 59016
rect 5448 58964 5500 59016
rect 9956 58896 10008 58948
rect 1400 58828 1452 58880
rect 2780 58828 2832 58880
rect 4213 58726 4265 58778
rect 4277 58726 4329 58778
rect 4341 58726 4393 58778
rect 4405 58726 4457 58778
rect 4469 58726 4521 58778
rect 7477 58726 7529 58778
rect 7541 58726 7593 58778
rect 7605 58726 7657 58778
rect 7669 58726 7721 58778
rect 7733 58726 7785 58778
rect 1768 58624 1820 58676
rect 1400 58488 1452 58540
rect 2228 58488 2280 58540
rect 4804 58488 4856 58540
rect 10140 58531 10192 58540
rect 10140 58497 10149 58531
rect 10149 58497 10183 58531
rect 10183 58497 10192 58531
rect 10140 58488 10192 58497
rect 1584 58284 1636 58336
rect 2504 58327 2556 58336
rect 2504 58293 2513 58327
rect 2513 58293 2547 58327
rect 2547 58293 2556 58327
rect 2504 58284 2556 58293
rect 2582 58182 2634 58234
rect 2646 58182 2698 58234
rect 2710 58182 2762 58234
rect 2774 58182 2826 58234
rect 2838 58182 2890 58234
rect 5845 58182 5897 58234
rect 5909 58182 5961 58234
rect 5973 58182 6025 58234
rect 6037 58182 6089 58234
rect 6101 58182 6153 58234
rect 9109 58182 9161 58234
rect 9173 58182 9225 58234
rect 9237 58182 9289 58234
rect 9301 58182 9353 58234
rect 9365 58182 9417 58234
rect 2136 58012 2188 58064
rect 2596 58012 2648 58064
rect 1492 57944 1544 57996
rect 1400 57919 1452 57928
rect 1400 57885 1409 57919
rect 1409 57885 1443 57919
rect 1443 57885 1452 57919
rect 1400 57876 1452 57885
rect 1676 57919 1728 57928
rect 1676 57885 1685 57919
rect 1685 57885 1719 57919
rect 1719 57885 1728 57919
rect 1676 57876 1728 57885
rect 2044 57944 2096 57996
rect 2320 57944 2372 57996
rect 2136 57808 2188 57860
rect 3516 57876 3568 57928
rect 2044 57740 2096 57792
rect 4213 57638 4265 57690
rect 4277 57638 4329 57690
rect 4341 57638 4393 57690
rect 4405 57638 4457 57690
rect 4469 57638 4521 57690
rect 7477 57638 7529 57690
rect 7541 57638 7593 57690
rect 7605 57638 7657 57690
rect 7669 57638 7721 57690
rect 7733 57638 7785 57690
rect 1400 57536 1452 57588
rect 2228 57536 2280 57588
rect 9864 57468 9916 57520
rect 1676 57443 1728 57452
rect 1676 57409 1685 57443
rect 1685 57409 1719 57443
rect 1719 57409 1728 57443
rect 1676 57400 1728 57409
rect 1492 57332 1544 57384
rect 2228 57400 2280 57452
rect 6184 57400 6236 57452
rect 10140 57443 10192 57452
rect 10140 57409 10149 57443
rect 10149 57409 10183 57443
rect 10183 57409 10192 57443
rect 10140 57400 10192 57409
rect 1400 57264 1452 57316
rect 3056 57332 3108 57384
rect 3148 57264 3200 57316
rect 3700 57196 3752 57248
rect 9956 57239 10008 57248
rect 9956 57205 9965 57239
rect 9965 57205 9999 57239
rect 9999 57205 10008 57239
rect 9956 57196 10008 57205
rect 2582 57094 2634 57146
rect 2646 57094 2698 57146
rect 2710 57094 2762 57146
rect 2774 57094 2826 57146
rect 2838 57094 2890 57146
rect 5845 57094 5897 57146
rect 5909 57094 5961 57146
rect 5973 57094 6025 57146
rect 6037 57094 6089 57146
rect 6101 57094 6153 57146
rect 9109 57094 9161 57146
rect 9173 57094 9225 57146
rect 9237 57094 9289 57146
rect 9301 57094 9353 57146
rect 9365 57094 9417 57146
rect 1676 56992 1728 57044
rect 1952 56992 2004 57044
rect 2136 56992 2188 57044
rect 9956 56992 10008 57044
rect 756 56856 808 56908
rect 1676 56856 1728 56908
rect 1492 56788 1544 56840
rect 1860 56788 1912 56840
rect 2228 56788 2280 56840
rect 6368 56788 6420 56840
rect 9956 56720 10008 56772
rect 664 56652 716 56704
rect 1308 56652 1360 56704
rect 1952 56652 2004 56704
rect 2504 56695 2556 56704
rect 2504 56661 2513 56695
rect 2513 56661 2547 56695
rect 2547 56661 2556 56695
rect 2504 56652 2556 56661
rect 3056 56652 3108 56704
rect 4712 56652 4764 56704
rect 4213 56550 4265 56602
rect 4277 56550 4329 56602
rect 4341 56550 4393 56602
rect 4405 56550 4457 56602
rect 4469 56550 4521 56602
rect 7477 56550 7529 56602
rect 7541 56550 7593 56602
rect 7605 56550 7657 56602
rect 7669 56550 7721 56602
rect 7733 56550 7785 56602
rect 1400 56448 1452 56500
rect 1860 56448 1912 56500
rect 3516 56448 3568 56500
rect 9956 56491 10008 56500
rect 9956 56457 9965 56491
rect 9965 56457 9999 56491
rect 9999 56457 10008 56491
rect 9956 56448 10008 56457
rect 1400 56312 1452 56364
rect 3148 56312 3200 56364
rect 10140 56355 10192 56364
rect 10140 56321 10149 56355
rect 10149 56321 10183 56355
rect 10183 56321 10192 56355
rect 10140 56312 10192 56321
rect 6552 56244 6604 56296
rect 2320 56219 2372 56228
rect 2320 56185 2329 56219
rect 2329 56185 2363 56219
rect 2363 56185 2372 56219
rect 2320 56176 2372 56185
rect 1492 56151 1544 56160
rect 1492 56117 1501 56151
rect 1501 56117 1535 56151
rect 1535 56117 1544 56151
rect 1492 56108 1544 56117
rect 2582 56006 2634 56058
rect 2646 56006 2698 56058
rect 2710 56006 2762 56058
rect 2774 56006 2826 56058
rect 2838 56006 2890 56058
rect 5845 56006 5897 56058
rect 5909 56006 5961 56058
rect 5973 56006 6025 56058
rect 6037 56006 6089 56058
rect 6101 56006 6153 56058
rect 9109 56006 9161 56058
rect 9173 56006 9225 56058
rect 9237 56006 9289 56058
rect 9301 56006 9353 56058
rect 9365 56006 9417 56058
rect 3056 55904 3108 55956
rect 3424 55904 3476 55956
rect 1492 55607 1544 55616
rect 1492 55573 1501 55607
rect 1501 55573 1535 55607
rect 1535 55573 1544 55607
rect 1492 55564 1544 55573
rect 3148 55564 3200 55616
rect 3700 55564 3752 55616
rect 4712 55564 4764 55616
rect 4213 55462 4265 55514
rect 4277 55462 4329 55514
rect 4341 55462 4393 55514
rect 4405 55462 4457 55514
rect 4469 55462 4521 55514
rect 7477 55462 7529 55514
rect 7541 55462 7593 55514
rect 7605 55462 7657 55514
rect 7669 55462 7721 55514
rect 7733 55462 7785 55514
rect 2964 55360 3016 55412
rect 3608 55360 3660 55412
rect 9864 55360 9916 55412
rect 7840 55292 7892 55344
rect 3148 55224 3200 55276
rect 10140 55267 10192 55276
rect 10140 55233 10149 55267
rect 10149 55233 10183 55267
rect 10183 55233 10192 55267
rect 10140 55224 10192 55233
rect 1492 55063 1544 55072
rect 1492 55029 1501 55063
rect 1501 55029 1535 55063
rect 1535 55029 1544 55063
rect 1492 55020 1544 55029
rect 2228 55063 2280 55072
rect 2228 55029 2237 55063
rect 2237 55029 2271 55063
rect 2271 55029 2280 55063
rect 2228 55020 2280 55029
rect 2582 54918 2634 54970
rect 2646 54918 2698 54970
rect 2710 54918 2762 54970
rect 2774 54918 2826 54970
rect 2838 54918 2890 54970
rect 5845 54918 5897 54970
rect 5909 54918 5961 54970
rect 5973 54918 6025 54970
rect 6037 54918 6089 54970
rect 6101 54918 6153 54970
rect 9109 54918 9161 54970
rect 9173 54918 9225 54970
rect 9237 54918 9289 54970
rect 9301 54918 9353 54970
rect 9365 54918 9417 54970
rect 3884 54816 3936 54868
rect 664 54612 716 54664
rect 3976 54612 4028 54664
rect 1400 54476 1452 54528
rect 4213 54374 4265 54426
rect 4277 54374 4329 54426
rect 4341 54374 4393 54426
rect 4405 54374 4457 54426
rect 4469 54374 4521 54426
rect 7477 54374 7529 54426
rect 7541 54374 7593 54426
rect 7605 54374 7657 54426
rect 7669 54374 7721 54426
rect 7733 54374 7785 54426
rect 7012 54136 7064 54188
rect 10140 54179 10192 54188
rect 10140 54145 10149 54179
rect 10149 54145 10183 54179
rect 10183 54145 10192 54179
rect 10140 54136 10192 54145
rect 7104 54068 7156 54120
rect 2228 54043 2280 54052
rect 2228 54009 2237 54043
rect 2237 54009 2271 54043
rect 2271 54009 2280 54043
rect 2228 54000 2280 54009
rect 1492 53975 1544 53984
rect 1492 53941 1501 53975
rect 1501 53941 1535 53975
rect 1535 53941 1544 53975
rect 1492 53932 1544 53941
rect 9956 53975 10008 53984
rect 9956 53941 9965 53975
rect 9965 53941 9999 53975
rect 9999 53941 10008 53975
rect 9956 53932 10008 53941
rect 2582 53830 2634 53882
rect 2646 53830 2698 53882
rect 2710 53830 2762 53882
rect 2774 53830 2826 53882
rect 2838 53830 2890 53882
rect 5845 53830 5897 53882
rect 5909 53830 5961 53882
rect 5973 53830 6025 53882
rect 6037 53830 6089 53882
rect 6101 53830 6153 53882
rect 9109 53830 9161 53882
rect 9173 53830 9225 53882
rect 9237 53830 9289 53882
rect 9301 53830 9353 53882
rect 9365 53830 9417 53882
rect 1216 53728 1268 53780
rect 1860 53728 1912 53780
rect 2044 53728 2096 53780
rect 2504 53728 2556 53780
rect 4068 53728 4120 53780
rect 2504 53592 2556 53644
rect 2964 53592 3016 53644
rect 2872 53567 2924 53576
rect 2872 53533 2881 53567
rect 2881 53533 2915 53567
rect 2915 53533 2924 53567
rect 2872 53524 2924 53533
rect 5448 53524 5500 53576
rect 7196 53456 7248 53508
rect 1400 53388 1452 53440
rect 2320 53431 2372 53440
rect 2320 53397 2329 53431
rect 2329 53397 2363 53431
rect 2363 53397 2372 53431
rect 2320 53388 2372 53397
rect 4213 53286 4265 53338
rect 4277 53286 4329 53338
rect 4341 53286 4393 53338
rect 4405 53286 4457 53338
rect 4469 53286 4521 53338
rect 7477 53286 7529 53338
rect 7541 53286 7593 53338
rect 7605 53286 7657 53338
rect 7669 53286 7721 53338
rect 7733 53286 7785 53338
rect 1952 53184 2004 53236
rect 3332 53184 3384 53236
rect 4068 53184 4120 53236
rect 5264 53184 5316 53236
rect 9956 53116 10008 53168
rect 1860 53048 1912 53100
rect 3056 53048 3108 53100
rect 3332 53091 3384 53100
rect 2044 52980 2096 53032
rect 3332 53057 3341 53091
rect 3341 53057 3375 53091
rect 3375 53057 3384 53091
rect 3332 53048 3384 53057
rect 4620 53048 4672 53100
rect 5264 53048 5316 53100
rect 10140 53091 10192 53100
rect 10140 53057 10149 53091
rect 10149 53057 10183 53091
rect 10183 53057 10192 53091
rect 10140 53048 10192 53057
rect 2872 52912 2924 52964
rect 2044 52844 2096 52896
rect 2964 52844 3016 52896
rect 5356 52912 5408 52964
rect 3332 52844 3384 52896
rect 9956 52887 10008 52896
rect 9956 52853 9965 52887
rect 9965 52853 9999 52887
rect 9999 52853 10008 52887
rect 9956 52844 10008 52853
rect 2582 52742 2634 52794
rect 2646 52742 2698 52794
rect 2710 52742 2762 52794
rect 2774 52742 2826 52794
rect 2838 52742 2890 52794
rect 5845 52742 5897 52794
rect 5909 52742 5961 52794
rect 5973 52742 6025 52794
rect 6037 52742 6089 52794
rect 6101 52742 6153 52794
rect 9109 52742 9161 52794
rect 9173 52742 9225 52794
rect 9237 52742 9289 52794
rect 9301 52742 9353 52794
rect 9365 52742 9417 52794
rect 3792 52683 3844 52692
rect 3792 52649 3801 52683
rect 3801 52649 3835 52683
rect 3835 52649 3844 52683
rect 3792 52640 3844 52649
rect 296 52572 348 52624
rect 1216 52572 1268 52624
rect 2596 52572 2648 52624
rect 2872 52572 2924 52624
rect 3884 52572 3936 52624
rect 5172 52572 5224 52624
rect 848 52436 900 52488
rect 1492 52436 1544 52488
rect 9956 52504 10008 52556
rect 1952 52479 2004 52488
rect 1952 52445 1961 52479
rect 1961 52445 1995 52479
rect 1995 52445 2004 52479
rect 1952 52436 2004 52445
rect 2596 52479 2648 52488
rect 2596 52445 2605 52479
rect 2605 52445 2639 52479
rect 2639 52445 2648 52479
rect 2596 52436 2648 52445
rect 3332 52436 3384 52488
rect 4620 52436 4672 52488
rect 2136 52368 2188 52420
rect 2320 52368 2372 52420
rect 4213 52198 4265 52250
rect 4277 52198 4329 52250
rect 4341 52198 4393 52250
rect 4405 52198 4457 52250
rect 4469 52198 4521 52250
rect 7477 52198 7529 52250
rect 7541 52198 7593 52250
rect 7605 52198 7657 52250
rect 7669 52198 7721 52250
rect 7733 52198 7785 52250
rect 2136 52096 2188 52148
rect 2412 51960 2464 52012
rect 10140 52003 10192 52012
rect 10140 51969 10149 52003
rect 10149 51969 10183 52003
rect 10183 51969 10192 52003
rect 10140 51960 10192 51969
rect 1492 51892 1544 51944
rect 1860 51892 1912 51944
rect 3332 51892 3384 51944
rect 3700 51824 3752 51876
rect 6644 51824 6696 51876
rect 1584 51756 1636 51808
rect 9956 51799 10008 51808
rect 9956 51765 9965 51799
rect 9965 51765 9999 51799
rect 9999 51765 10008 51799
rect 9956 51756 10008 51765
rect 2582 51654 2634 51706
rect 2646 51654 2698 51706
rect 2710 51654 2762 51706
rect 2774 51654 2826 51706
rect 2838 51654 2890 51706
rect 5845 51654 5897 51706
rect 5909 51654 5961 51706
rect 5973 51654 6025 51706
rect 6037 51654 6089 51706
rect 6101 51654 6153 51706
rect 9109 51654 9161 51706
rect 9173 51654 9225 51706
rect 9237 51654 9289 51706
rect 9301 51654 9353 51706
rect 9365 51654 9417 51706
rect 1952 51552 2004 51604
rect 3792 51552 3844 51604
rect 9864 51552 9916 51604
rect 1584 51391 1636 51400
rect 1584 51357 1593 51391
rect 1593 51357 1627 51391
rect 1627 51357 1636 51391
rect 1584 51348 1636 51357
rect 1768 51391 1820 51400
rect 1768 51357 1777 51391
rect 1777 51357 1811 51391
rect 1811 51357 1820 51391
rect 1768 51348 1820 51357
rect 3700 51484 3752 51536
rect 3976 51484 4028 51536
rect 5540 51484 5592 51536
rect 5816 51484 5868 51536
rect 3792 51391 3844 51400
rect 3792 51357 3801 51391
rect 3801 51357 3835 51391
rect 3835 51357 3844 51391
rect 3792 51348 3844 51357
rect 1676 51323 1728 51332
rect 1676 51289 1685 51323
rect 1685 51289 1719 51323
rect 1719 51289 1728 51323
rect 1676 51280 1728 51289
rect 2320 51280 2372 51332
rect 9956 51280 10008 51332
rect 2136 51212 2188 51264
rect 2596 51212 2648 51264
rect 3976 51255 4028 51264
rect 3976 51221 3985 51255
rect 3985 51221 4019 51255
rect 4019 51221 4028 51255
rect 3976 51212 4028 51221
rect 4213 51110 4265 51162
rect 4277 51110 4329 51162
rect 4341 51110 4393 51162
rect 4405 51110 4457 51162
rect 4469 51110 4521 51162
rect 7477 51110 7529 51162
rect 7541 51110 7593 51162
rect 7605 51110 7657 51162
rect 7669 51110 7721 51162
rect 7733 51110 7785 51162
rect 1308 51008 1360 51060
rect 3424 51051 3476 51060
rect 3424 51017 3433 51051
rect 3433 51017 3467 51051
rect 3467 51017 3476 51051
rect 3424 51008 3476 51017
rect 9864 51008 9916 51060
rect 2964 50872 3016 50924
rect 1860 50804 1912 50856
rect 1676 50736 1728 50788
rect 2596 50736 2648 50788
rect 3056 50736 3108 50788
rect 3884 50804 3936 50856
rect 5172 50872 5224 50924
rect 5540 50872 5592 50924
rect 10140 50915 10192 50924
rect 10140 50881 10149 50915
rect 10149 50881 10183 50915
rect 10183 50881 10192 50915
rect 10140 50872 10192 50881
rect 4160 50736 4212 50788
rect 5448 50668 5500 50720
rect 5816 50736 5868 50788
rect 6736 50736 6788 50788
rect 2582 50566 2634 50618
rect 2646 50566 2698 50618
rect 2710 50566 2762 50618
rect 2774 50566 2826 50618
rect 2838 50566 2890 50618
rect 5845 50566 5897 50618
rect 5909 50566 5961 50618
rect 5973 50566 6025 50618
rect 6037 50566 6089 50618
rect 6101 50566 6153 50618
rect 9109 50566 9161 50618
rect 9173 50566 9225 50618
rect 9237 50566 9289 50618
rect 9301 50566 9353 50618
rect 9365 50566 9417 50618
rect 1768 50328 1820 50380
rect 3332 50328 3384 50380
rect 3792 50371 3844 50380
rect 3792 50337 3801 50371
rect 3801 50337 3835 50371
rect 3835 50337 3844 50371
rect 3792 50328 3844 50337
rect 3884 50328 3936 50380
rect 1860 50260 1912 50312
rect 2596 50260 2648 50312
rect 3240 50260 3292 50312
rect 4160 50260 4212 50312
rect 1216 50124 1268 50176
rect 9956 50192 10008 50244
rect 1952 50124 2004 50176
rect 2504 50167 2556 50176
rect 2504 50133 2513 50167
rect 2513 50133 2547 50167
rect 2547 50133 2556 50167
rect 2504 50124 2556 50133
rect 4213 50022 4265 50074
rect 4277 50022 4329 50074
rect 4341 50022 4393 50074
rect 4405 50022 4457 50074
rect 4469 50022 4521 50074
rect 7477 50022 7529 50074
rect 7541 50022 7593 50074
rect 7605 50022 7657 50074
rect 7669 50022 7721 50074
rect 7733 50022 7785 50074
rect 1492 49963 1544 49972
rect 1492 49929 1501 49963
rect 1501 49929 1535 49963
rect 1535 49929 1544 49963
rect 1492 49920 1544 49929
rect 3700 49920 3752 49972
rect 9956 49963 10008 49972
rect 9956 49929 9965 49963
rect 9965 49929 9999 49963
rect 9999 49929 10008 49963
rect 9956 49920 10008 49929
rect 1952 49716 2004 49768
rect 2228 49716 2280 49768
rect 2688 49784 2740 49836
rect 2964 49784 3016 49836
rect 3424 49716 3476 49768
rect 6460 49784 6512 49836
rect 3884 49716 3936 49768
rect 204 49648 256 49700
rect 2688 49648 2740 49700
rect 2872 49648 2924 49700
rect 3700 49648 3752 49700
rect 10140 49648 10192 49700
rect 2228 49623 2280 49632
rect 2228 49589 2237 49623
rect 2237 49589 2271 49623
rect 2271 49589 2280 49623
rect 2228 49580 2280 49589
rect 2582 49478 2634 49530
rect 2646 49478 2698 49530
rect 2710 49478 2762 49530
rect 2774 49478 2826 49530
rect 2838 49478 2890 49530
rect 5845 49478 5897 49530
rect 5909 49478 5961 49530
rect 5973 49478 6025 49530
rect 6037 49478 6089 49530
rect 6101 49478 6153 49530
rect 9109 49478 9161 49530
rect 9173 49478 9225 49530
rect 9237 49478 9289 49530
rect 9301 49478 9353 49530
rect 9365 49478 9417 49530
rect 1400 49376 1452 49428
rect 1860 49376 1912 49428
rect 3240 49376 3292 49428
rect 1124 49240 1176 49292
rect 1400 49240 1452 49292
rect 2780 49240 2832 49292
rect 3792 49283 3844 49292
rect 3792 49249 3801 49283
rect 3801 49249 3835 49283
rect 3835 49249 3844 49283
rect 3792 49240 3844 49249
rect 1124 49104 1176 49156
rect 2964 49172 3016 49224
rect 1492 49079 1544 49088
rect 1492 49045 1501 49079
rect 1501 49045 1535 49079
rect 1535 49045 1544 49079
rect 1492 49036 1544 49045
rect 2872 49104 2924 49156
rect 3884 49172 3936 49224
rect 4213 48934 4265 48986
rect 4277 48934 4329 48986
rect 4341 48934 4393 48986
rect 4405 48934 4457 48986
rect 4469 48934 4521 48986
rect 7477 48934 7529 48986
rect 7541 48934 7593 48986
rect 7605 48934 7657 48986
rect 7669 48934 7721 48986
rect 7733 48934 7785 48986
rect 2780 48764 2832 48816
rect 4528 48764 4580 48816
rect 3700 48696 3752 48748
rect 10140 48739 10192 48748
rect 10140 48705 10149 48739
rect 10149 48705 10183 48739
rect 10183 48705 10192 48739
rect 10140 48696 10192 48705
rect 6828 48628 6880 48680
rect 2228 48603 2280 48612
rect 2228 48569 2237 48603
rect 2237 48569 2271 48603
rect 2271 48569 2280 48603
rect 2228 48560 2280 48569
rect 1492 48535 1544 48544
rect 1492 48501 1501 48535
rect 1501 48501 1535 48535
rect 1535 48501 1544 48535
rect 1492 48492 1544 48501
rect 2582 48390 2634 48442
rect 2646 48390 2698 48442
rect 2710 48390 2762 48442
rect 2774 48390 2826 48442
rect 2838 48390 2890 48442
rect 5845 48390 5897 48442
rect 5909 48390 5961 48442
rect 5973 48390 6025 48442
rect 6037 48390 6089 48442
rect 6101 48390 6153 48442
rect 9109 48390 9161 48442
rect 9173 48390 9225 48442
rect 9237 48390 9289 48442
rect 9301 48390 9353 48442
rect 9365 48390 9417 48442
rect 1768 48288 1820 48340
rect 2504 48263 2556 48272
rect 2504 48229 2513 48263
rect 2513 48229 2547 48263
rect 2547 48229 2556 48263
rect 2504 48220 2556 48229
rect 756 48152 808 48204
rect 1676 48127 1728 48136
rect 1676 48093 1685 48127
rect 1685 48093 1719 48127
rect 1719 48093 1728 48127
rect 1676 48084 1728 48093
rect 2872 48016 2924 48068
rect 1492 47991 1544 48000
rect 1492 47957 1501 47991
rect 1501 47957 1535 47991
rect 1535 47957 1544 47991
rect 1492 47948 1544 47957
rect 2780 47948 2832 48000
rect 3332 47948 3384 48000
rect 4213 47846 4265 47898
rect 4277 47846 4329 47898
rect 4341 47846 4393 47898
rect 4405 47846 4457 47898
rect 4469 47846 4521 47898
rect 7477 47846 7529 47898
rect 7541 47846 7593 47898
rect 7605 47846 7657 47898
rect 7669 47846 7721 47898
rect 7733 47846 7785 47898
rect 664 47744 716 47796
rect 3332 47744 3384 47796
rect 2964 47719 3016 47728
rect 2964 47685 2973 47719
rect 2973 47685 3007 47719
rect 3007 47685 3016 47719
rect 2964 47676 3016 47685
rect 1400 47608 1452 47660
rect 2780 47608 2832 47660
rect 2872 47651 2924 47660
rect 2872 47617 2881 47651
rect 2881 47617 2915 47651
rect 2915 47617 2924 47651
rect 2872 47608 2924 47617
rect 10140 47651 10192 47660
rect 848 47472 900 47524
rect 10140 47617 10149 47651
rect 10149 47617 10183 47651
rect 10183 47617 10192 47651
rect 10140 47608 10192 47617
rect 1492 47447 1544 47456
rect 1492 47413 1501 47447
rect 1501 47413 1535 47447
rect 1535 47413 1544 47447
rect 1492 47404 1544 47413
rect 2228 47447 2280 47456
rect 2228 47413 2237 47447
rect 2237 47413 2271 47447
rect 2271 47413 2280 47447
rect 2228 47404 2280 47413
rect 2582 47302 2634 47354
rect 2646 47302 2698 47354
rect 2710 47302 2762 47354
rect 2774 47302 2826 47354
rect 2838 47302 2890 47354
rect 5845 47302 5897 47354
rect 5909 47302 5961 47354
rect 5973 47302 6025 47354
rect 6037 47302 6089 47354
rect 6101 47302 6153 47354
rect 9109 47302 9161 47354
rect 9173 47302 9225 47354
rect 9237 47302 9289 47354
rect 9301 47302 9353 47354
rect 9365 47302 9417 47354
rect 1676 47200 1728 47252
rect 3424 47200 3476 47252
rect 1032 47064 1084 47116
rect 1584 46996 1636 47048
rect 4896 47132 4948 47184
rect 3884 46996 3936 47048
rect 204 46767 256 46776
rect 204 46733 213 46767
rect 213 46733 247 46767
rect 247 46733 256 46767
rect 204 46724 256 46733
rect 2964 46928 3016 46980
rect 1308 46860 1360 46912
rect 2780 46860 2832 46912
rect 8300 46860 8352 46912
rect 4213 46758 4265 46810
rect 4277 46758 4329 46810
rect 4341 46758 4393 46810
rect 4405 46758 4457 46810
rect 4469 46758 4521 46810
rect 7477 46758 7529 46810
rect 7541 46758 7593 46810
rect 7605 46758 7657 46810
rect 7669 46758 7721 46810
rect 7733 46758 7785 46810
rect 1124 46656 1176 46708
rect 3700 46699 3752 46708
rect 3700 46665 3709 46699
rect 3709 46665 3743 46699
rect 3743 46665 3752 46699
rect 3700 46656 3752 46665
rect 204 46588 256 46640
rect 2780 46520 2832 46572
rect 3056 46520 3108 46572
rect 3884 46588 3936 46640
rect 10140 46563 10192 46572
rect 10140 46529 10149 46563
rect 10149 46529 10183 46563
rect 10183 46529 10192 46563
rect 10140 46520 10192 46529
rect 3056 46427 3108 46436
rect 1400 46316 1452 46368
rect 2228 46359 2280 46368
rect 2228 46325 2237 46359
rect 2237 46325 2271 46359
rect 2271 46325 2280 46359
rect 2228 46316 2280 46325
rect 3056 46393 3065 46427
rect 3065 46393 3099 46427
rect 3099 46393 3108 46427
rect 3056 46384 3108 46393
rect 6736 46384 6788 46436
rect 4620 46316 4672 46368
rect 4896 46316 4948 46368
rect 9956 46359 10008 46368
rect 9956 46325 9965 46359
rect 9965 46325 9999 46359
rect 9999 46325 10008 46359
rect 9956 46316 10008 46325
rect 296 46180 348 46232
rect 664 46180 716 46232
rect 2582 46214 2634 46266
rect 2646 46214 2698 46266
rect 2710 46214 2762 46266
rect 2774 46214 2826 46266
rect 2838 46214 2890 46266
rect 5845 46214 5897 46266
rect 5909 46214 5961 46266
rect 5973 46214 6025 46266
rect 6037 46214 6089 46266
rect 6101 46214 6153 46266
rect 9109 46214 9161 46266
rect 9173 46214 9225 46266
rect 9237 46214 9289 46266
rect 9301 46214 9353 46266
rect 9365 46214 9417 46266
rect 112 46112 164 46164
rect 3056 46112 3108 46164
rect 3240 46112 3292 46164
rect 4620 46112 4672 46164
rect 5080 46112 5132 46164
rect 296 46044 348 46096
rect 2412 46019 2464 46028
rect 2412 45985 2421 46019
rect 2421 45985 2455 46019
rect 2455 45985 2464 46019
rect 2412 45976 2464 45985
rect 3332 45976 3384 46028
rect 3516 45976 3568 46028
rect 1584 45908 1636 45960
rect 1492 45815 1544 45824
rect 1492 45781 1501 45815
rect 1501 45781 1535 45815
rect 1535 45781 1544 45815
rect 1492 45772 1544 45781
rect 2228 45772 2280 45824
rect 3148 45908 3200 45960
rect 3240 45908 3292 45960
rect 3700 45908 3752 45960
rect 4213 45670 4265 45722
rect 4277 45670 4329 45722
rect 4341 45670 4393 45722
rect 4405 45670 4457 45722
rect 4469 45670 4521 45722
rect 7477 45670 7529 45722
rect 7541 45670 7593 45722
rect 7605 45670 7657 45722
rect 7669 45670 7721 45722
rect 7733 45670 7785 45722
rect 388 45568 440 45620
rect 1584 45568 1636 45620
rect 3332 45500 3384 45552
rect 5540 45500 5592 45552
rect 3976 45432 4028 45484
rect 10140 45475 10192 45484
rect 10140 45441 10149 45475
rect 10149 45441 10183 45475
rect 10183 45441 10192 45475
rect 10140 45432 10192 45441
rect 2412 45407 2464 45416
rect 2412 45373 2421 45407
rect 2421 45373 2455 45407
rect 2455 45373 2464 45407
rect 2412 45364 2464 45373
rect 9864 45228 9916 45280
rect 2582 45126 2634 45178
rect 2646 45126 2698 45178
rect 2710 45126 2762 45178
rect 2774 45126 2826 45178
rect 2838 45126 2890 45178
rect 5845 45126 5897 45178
rect 5909 45126 5961 45178
rect 5973 45126 6025 45178
rect 6037 45126 6089 45178
rect 6101 45126 6153 45178
rect 9109 45126 9161 45178
rect 9173 45126 9225 45178
rect 9237 45126 9289 45178
rect 9301 45126 9353 45178
rect 9365 45126 9417 45178
rect 1308 45024 1360 45076
rect 2964 45024 3016 45076
rect 2228 44888 2280 44940
rect 2596 44888 2648 44940
rect 2412 44820 2464 44872
rect 3792 44820 3844 44872
rect 1400 44727 1452 44736
rect 1400 44693 1409 44727
rect 1409 44693 1443 44727
rect 1443 44693 1452 44727
rect 1400 44684 1452 44693
rect 1584 44684 1636 44736
rect 4213 44582 4265 44634
rect 4277 44582 4329 44634
rect 4341 44582 4393 44634
rect 4405 44582 4457 44634
rect 4469 44582 4521 44634
rect 7477 44582 7529 44634
rect 7541 44582 7593 44634
rect 7605 44582 7657 44634
rect 7669 44582 7721 44634
rect 7733 44582 7785 44634
rect 112 44412 164 44464
rect 848 44412 900 44464
rect 2596 44480 2648 44532
rect 1676 44455 1728 44464
rect 1676 44421 1685 44455
rect 1685 44421 1719 44455
rect 1719 44421 1728 44455
rect 1676 44412 1728 44421
rect 2504 44412 2556 44464
rect 1492 44344 1544 44396
rect 2412 44344 2464 44396
rect 2596 44387 2648 44396
rect 2596 44353 2605 44387
rect 2605 44353 2639 44387
rect 2639 44353 2648 44387
rect 2596 44344 2648 44353
rect 9956 44412 10008 44464
rect 10140 44387 10192 44396
rect 2504 44208 2556 44260
rect 10140 44353 10149 44387
rect 10149 44353 10183 44387
rect 10183 44353 10192 44387
rect 10140 44344 10192 44353
rect 1860 44140 1912 44192
rect 2412 44183 2464 44192
rect 2412 44149 2421 44183
rect 2421 44149 2455 44183
rect 2455 44149 2464 44183
rect 2412 44140 2464 44149
rect 9956 44183 10008 44192
rect 9956 44149 9965 44183
rect 9965 44149 9999 44183
rect 9999 44149 10008 44183
rect 9956 44140 10008 44149
rect 2582 44038 2634 44090
rect 2646 44038 2698 44090
rect 2710 44038 2762 44090
rect 2774 44038 2826 44090
rect 2838 44038 2890 44090
rect 5845 44038 5897 44090
rect 5909 44038 5961 44090
rect 5973 44038 6025 44090
rect 6037 44038 6089 44090
rect 6101 44038 6153 44090
rect 9109 44038 9161 44090
rect 9173 44038 9225 44090
rect 9237 44038 9289 44090
rect 9301 44038 9353 44090
rect 9365 44038 9417 44090
rect 1492 43732 1544 43784
rect 1676 43775 1728 43784
rect 1676 43741 1685 43775
rect 1685 43741 1719 43775
rect 1719 43741 1728 43775
rect 2504 43800 2556 43852
rect 1676 43732 1728 43741
rect 2228 43732 2280 43784
rect 4068 43732 4120 43784
rect 9956 43664 10008 43716
rect 1584 43596 1636 43648
rect 2780 43596 2832 43648
rect 3976 43639 4028 43648
rect 3976 43605 3985 43639
rect 3985 43605 4019 43639
rect 4019 43605 4028 43639
rect 3976 43596 4028 43605
rect 4213 43494 4265 43546
rect 4277 43494 4329 43546
rect 4341 43494 4393 43546
rect 4405 43494 4457 43546
rect 4469 43494 4521 43546
rect 7477 43494 7529 43546
rect 7541 43494 7593 43546
rect 7605 43494 7657 43546
rect 7669 43494 7721 43546
rect 7733 43494 7785 43546
rect 9864 43392 9916 43444
rect 4160 43324 4212 43376
rect 4988 43324 5040 43376
rect 1492 43256 1544 43308
rect 2504 43256 2556 43308
rect 3148 43256 3200 43308
rect 9864 43299 9916 43308
rect 9864 43265 9873 43299
rect 9873 43265 9907 43299
rect 9907 43265 9916 43299
rect 9864 43256 9916 43265
rect 8484 43188 8536 43240
rect 2504 43095 2556 43104
rect 2504 43061 2513 43095
rect 2513 43061 2547 43095
rect 2547 43061 2556 43095
rect 2504 43052 2556 43061
rect 10048 43095 10100 43104
rect 10048 43061 10057 43095
rect 10057 43061 10091 43095
rect 10091 43061 10100 43095
rect 10048 43052 10100 43061
rect 2582 42950 2634 43002
rect 2646 42950 2698 43002
rect 2710 42950 2762 43002
rect 2774 42950 2826 43002
rect 2838 42950 2890 43002
rect 5845 42950 5897 43002
rect 5909 42950 5961 43002
rect 5973 42950 6025 43002
rect 6037 42950 6089 43002
rect 6101 42950 6153 43002
rect 9109 42950 9161 43002
rect 9173 42950 9225 43002
rect 9237 42950 9289 43002
rect 9301 42950 9353 43002
rect 9365 42950 9417 43002
rect 20 42780 72 42832
rect 940 42712 992 42764
rect 20 42644 72 42696
rect 756 42644 808 42696
rect 940 42440 992 42492
rect 296 42372 348 42424
rect 848 42372 900 42424
rect 1676 42687 1728 42696
rect 1676 42653 1685 42687
rect 1685 42653 1719 42687
rect 1719 42653 1728 42687
rect 1676 42644 1728 42653
rect 4988 42644 5040 42696
rect 9864 42712 9916 42764
rect 8392 42644 8444 42696
rect 5448 42576 5500 42628
rect 1492 42551 1544 42560
rect 1492 42517 1501 42551
rect 1501 42517 1535 42551
rect 1535 42517 1544 42551
rect 1492 42508 1544 42517
rect 2228 42551 2280 42560
rect 2228 42517 2237 42551
rect 2237 42517 2271 42551
rect 2271 42517 2280 42551
rect 2228 42508 2280 42517
rect 4213 42406 4265 42458
rect 4277 42406 4329 42458
rect 4341 42406 4393 42458
rect 4405 42406 4457 42458
rect 4469 42406 4521 42458
rect 7477 42406 7529 42458
rect 7541 42406 7593 42458
rect 7605 42406 7657 42458
rect 7669 42406 7721 42458
rect 7733 42406 7785 42458
rect 1676 42304 1728 42356
rect 6920 42304 6972 42356
rect 4896 42236 4948 42288
rect 5080 42236 5132 42288
rect 4988 42168 5040 42220
rect 1400 42100 1452 42152
rect 1584 42100 1636 42152
rect 1400 41964 1452 42016
rect 10048 42007 10100 42016
rect 10048 41973 10057 42007
rect 10057 41973 10091 42007
rect 10091 41973 10100 42007
rect 10048 41964 10100 41973
rect 2582 41862 2634 41914
rect 2646 41862 2698 41914
rect 2710 41862 2762 41914
rect 2774 41862 2826 41914
rect 2838 41862 2890 41914
rect 5845 41862 5897 41914
rect 5909 41862 5961 41914
rect 5973 41862 6025 41914
rect 6037 41862 6089 41914
rect 6101 41862 6153 41914
rect 9109 41862 9161 41914
rect 9173 41862 9225 41914
rect 9237 41862 9289 41914
rect 9301 41862 9353 41914
rect 9365 41862 9417 41914
rect 1952 41692 2004 41744
rect 2320 41692 2372 41744
rect 6736 41556 6788 41608
rect 1216 41488 1268 41540
rect 1952 41488 2004 41540
rect 3792 41488 3844 41540
rect 5264 41488 5316 41540
rect 1492 41463 1544 41472
rect 1492 41429 1501 41463
rect 1501 41429 1535 41463
rect 1535 41429 1544 41463
rect 1492 41420 1544 41429
rect 4213 41318 4265 41370
rect 4277 41318 4329 41370
rect 4341 41318 4393 41370
rect 4405 41318 4457 41370
rect 4469 41318 4521 41370
rect 7477 41318 7529 41370
rect 7541 41318 7593 41370
rect 7605 41318 7657 41370
rect 7669 41318 7721 41370
rect 7733 41318 7785 41370
rect 8576 41216 8628 41268
rect 4896 41148 4948 41200
rect 5356 41148 5408 41200
rect 4988 41080 5040 41132
rect 1492 40919 1544 40928
rect 1492 40885 1501 40919
rect 1501 40885 1535 40919
rect 1535 40885 1544 40919
rect 1492 40876 1544 40885
rect 10048 40919 10100 40928
rect 10048 40885 10057 40919
rect 10057 40885 10091 40919
rect 10091 40885 10100 40919
rect 10048 40876 10100 40885
rect 2582 40774 2634 40826
rect 2646 40774 2698 40826
rect 2710 40774 2762 40826
rect 2774 40774 2826 40826
rect 2838 40774 2890 40826
rect 5845 40774 5897 40826
rect 5909 40774 5961 40826
rect 5973 40774 6025 40826
rect 6037 40774 6089 40826
rect 6101 40774 6153 40826
rect 9109 40774 9161 40826
rect 9173 40774 9225 40826
rect 9237 40774 9289 40826
rect 9301 40774 9353 40826
rect 9365 40774 9417 40826
rect 112 40672 164 40724
rect 1308 40672 1360 40724
rect 3424 40672 3476 40724
rect 3976 40672 4028 40724
rect 4804 40672 4856 40724
rect 5356 40672 5408 40724
rect 296 40604 348 40656
rect 1124 40604 1176 40656
rect 1032 40536 1084 40588
rect 1400 40536 1452 40588
rect 8668 40468 8720 40520
rect 1400 40400 1452 40452
rect 2504 40400 2556 40452
rect 1492 40375 1544 40384
rect 1492 40341 1501 40375
rect 1501 40341 1535 40375
rect 1535 40341 1544 40375
rect 1492 40332 1544 40341
rect 2412 40332 2464 40384
rect 3792 40332 3844 40384
rect 4213 40230 4265 40282
rect 4277 40230 4329 40282
rect 4341 40230 4393 40282
rect 4405 40230 4457 40282
rect 4469 40230 4521 40282
rect 7477 40230 7529 40282
rect 7541 40230 7593 40282
rect 7605 40230 7657 40282
rect 7669 40230 7721 40282
rect 7733 40230 7785 40282
rect 1676 40128 1728 40180
rect 1860 40128 1912 40180
rect 4620 40128 4672 40180
rect 2412 40060 2464 40112
rect 2504 40035 2556 40044
rect 2504 40001 2513 40035
rect 2513 40001 2547 40035
rect 2547 40001 2556 40035
rect 2504 39992 2556 40001
rect 4804 40060 4856 40112
rect 1492 39831 1544 39840
rect 1492 39797 1501 39831
rect 1501 39797 1535 39831
rect 1535 39797 1544 39831
rect 1492 39788 1544 39797
rect 2582 39686 2634 39738
rect 2646 39686 2698 39738
rect 2710 39686 2762 39738
rect 2774 39686 2826 39738
rect 2838 39686 2890 39738
rect 5845 39686 5897 39738
rect 5909 39686 5961 39738
rect 5973 39686 6025 39738
rect 6037 39686 6089 39738
rect 6101 39686 6153 39738
rect 9109 39686 9161 39738
rect 9173 39686 9225 39738
rect 9237 39686 9289 39738
rect 9301 39686 9353 39738
rect 9365 39686 9417 39738
rect 5724 39516 5776 39568
rect 3240 39448 3292 39500
rect 2504 39423 2556 39432
rect 2504 39389 2513 39423
rect 2513 39389 2547 39423
rect 2547 39389 2556 39423
rect 2504 39380 2556 39389
rect 2964 39380 3016 39432
rect 9864 39423 9916 39432
rect 9864 39389 9873 39423
rect 9873 39389 9907 39423
rect 9907 39389 9916 39423
rect 9864 39380 9916 39389
rect 1492 39287 1544 39296
rect 1492 39253 1501 39287
rect 1501 39253 1535 39287
rect 1535 39253 1544 39287
rect 1492 39244 1544 39253
rect 10048 39287 10100 39296
rect 10048 39253 10057 39287
rect 10057 39253 10091 39287
rect 10091 39253 10100 39287
rect 10048 39244 10100 39253
rect 4213 39142 4265 39194
rect 4277 39142 4329 39194
rect 4341 39142 4393 39194
rect 4405 39142 4457 39194
rect 4469 39142 4521 39194
rect 7477 39142 7529 39194
rect 7541 39142 7593 39194
rect 7605 39142 7657 39194
rect 7669 39142 7721 39194
rect 7733 39142 7785 39194
rect 940 38972 992 39024
rect 2412 38972 2464 39024
rect 1584 38904 1636 38956
rect 2504 38947 2556 38956
rect 2504 38913 2513 38947
rect 2513 38913 2547 38947
rect 2547 38913 2556 38947
rect 2504 38904 2556 38913
rect 4620 38904 4672 38956
rect 4804 38836 4856 38888
rect 1492 38811 1544 38820
rect 1492 38777 1501 38811
rect 1501 38777 1535 38811
rect 1535 38777 1544 38811
rect 1492 38768 1544 38777
rect 2964 38700 3016 38752
rect 4252 38700 4304 38752
rect 9864 38700 9916 38752
rect 2582 38598 2634 38650
rect 2646 38598 2698 38650
rect 2710 38598 2762 38650
rect 2774 38598 2826 38650
rect 2838 38598 2890 38650
rect 5845 38598 5897 38650
rect 5909 38598 5961 38650
rect 5973 38598 6025 38650
rect 6037 38598 6089 38650
rect 6101 38598 6153 38650
rect 9109 38598 9161 38650
rect 9173 38598 9225 38650
rect 9237 38598 9289 38650
rect 9301 38598 9353 38650
rect 9365 38598 9417 38650
rect 7380 38428 7432 38480
rect 2228 38360 2280 38412
rect 2504 38335 2556 38344
rect 2504 38301 2513 38335
rect 2513 38301 2547 38335
rect 2547 38301 2556 38335
rect 2504 38292 2556 38301
rect 4252 38335 4304 38344
rect 2228 38224 2280 38276
rect 4252 38301 4261 38335
rect 4261 38301 4295 38335
rect 4295 38301 4304 38335
rect 4252 38292 4304 38301
rect 4620 38292 4672 38344
rect 1492 38199 1544 38208
rect 1492 38165 1501 38199
rect 1501 38165 1535 38199
rect 1535 38165 1544 38199
rect 1492 38156 1544 38165
rect 10048 38199 10100 38208
rect 10048 38165 10057 38199
rect 10057 38165 10091 38199
rect 10091 38165 10100 38199
rect 10048 38156 10100 38165
rect 4213 38054 4265 38106
rect 4277 38054 4329 38106
rect 4341 38054 4393 38106
rect 4405 38054 4457 38106
rect 4469 38054 4521 38106
rect 7477 38054 7529 38106
rect 7541 38054 7593 38106
rect 7605 38054 7657 38106
rect 7669 38054 7721 38106
rect 7733 38054 7785 38106
rect 1400 37952 1452 38004
rect 4068 37952 4120 38004
rect 1860 37884 1912 37936
rect 2320 37884 2372 37936
rect 2504 37859 2556 37868
rect 1492 37748 1544 37800
rect 1860 37748 1912 37800
rect 2504 37825 2513 37859
rect 2513 37825 2547 37859
rect 2547 37825 2556 37859
rect 2504 37816 2556 37825
rect 3700 37816 3752 37868
rect 4160 37859 4212 37868
rect 4160 37825 4169 37859
rect 4169 37825 4203 37859
rect 4203 37825 4212 37859
rect 4160 37816 4212 37825
rect 4620 37816 4672 37868
rect 3240 37655 3292 37664
rect 3240 37621 3249 37655
rect 3249 37621 3283 37655
rect 3283 37621 3292 37655
rect 3240 37612 3292 37621
rect 9864 37612 9916 37664
rect 2582 37510 2634 37562
rect 2646 37510 2698 37562
rect 2710 37510 2762 37562
rect 2774 37510 2826 37562
rect 2838 37510 2890 37562
rect 5845 37510 5897 37562
rect 5909 37510 5961 37562
rect 5973 37510 6025 37562
rect 6037 37510 6089 37562
rect 6101 37510 6153 37562
rect 9109 37510 9161 37562
rect 9173 37510 9225 37562
rect 9237 37510 9289 37562
rect 9301 37510 9353 37562
rect 9365 37510 9417 37562
rect 1492 37272 1544 37324
rect 2044 37204 2096 37256
rect 2964 37247 3016 37256
rect 2964 37213 2973 37247
rect 2973 37213 3007 37247
rect 3007 37213 3016 37247
rect 2964 37204 3016 37213
rect 3792 37204 3844 37256
rect 9864 37247 9916 37256
rect 9864 37213 9873 37247
rect 9873 37213 9907 37247
rect 9907 37213 9916 37247
rect 9864 37204 9916 37213
rect 2412 37136 2464 37188
rect 4160 37136 4212 37188
rect 1584 37111 1636 37120
rect 1584 37077 1593 37111
rect 1593 37077 1627 37111
rect 1627 37077 1636 37111
rect 1584 37068 1636 37077
rect 2320 37111 2372 37120
rect 2320 37077 2329 37111
rect 2329 37077 2363 37111
rect 2363 37077 2372 37111
rect 2320 37068 2372 37077
rect 2964 37068 3016 37120
rect 3148 37068 3200 37120
rect 10048 37111 10100 37120
rect 10048 37077 10057 37111
rect 10057 37077 10091 37111
rect 10091 37077 10100 37111
rect 10048 37068 10100 37077
rect 4213 36966 4265 37018
rect 4277 36966 4329 37018
rect 4341 36966 4393 37018
rect 4405 36966 4457 37018
rect 4469 36966 4521 37018
rect 7477 36966 7529 37018
rect 7541 36966 7593 37018
rect 7605 36966 7657 37018
rect 7669 36966 7721 37018
rect 7733 36966 7785 37018
rect 2412 36864 2464 36916
rect 4804 36864 4856 36916
rect 1768 36728 1820 36780
rect 2044 36728 2096 36780
rect 2412 36728 2464 36780
rect 3516 36728 3568 36780
rect 2228 36660 2280 36712
rect 4620 36728 4672 36780
rect 1492 36567 1544 36576
rect 1492 36533 1501 36567
rect 1501 36533 1535 36567
rect 1535 36533 1544 36567
rect 1492 36524 1544 36533
rect 1676 36524 1728 36576
rect 1860 36524 1912 36576
rect 9864 36524 9916 36576
rect 2582 36422 2634 36474
rect 2646 36422 2698 36474
rect 2710 36422 2762 36474
rect 2774 36422 2826 36474
rect 2838 36422 2890 36474
rect 5845 36422 5897 36474
rect 5909 36422 5961 36474
rect 5973 36422 6025 36474
rect 6037 36422 6089 36474
rect 6101 36422 6153 36474
rect 9109 36422 9161 36474
rect 9173 36422 9225 36474
rect 9237 36422 9289 36474
rect 9301 36422 9353 36474
rect 9365 36422 9417 36474
rect 1400 36320 1452 36372
rect 1676 36320 1728 36372
rect 2228 36363 2280 36372
rect 2228 36329 2237 36363
rect 2237 36329 2271 36363
rect 2271 36329 2280 36363
rect 2228 36320 2280 36329
rect 1952 36116 2004 36168
rect 2228 36116 2280 36168
rect 1584 36023 1636 36032
rect 1584 35989 1593 36023
rect 1593 35989 1627 36023
rect 1627 35989 1636 36023
rect 1584 35980 1636 35989
rect 1768 36048 1820 36100
rect 4620 36116 4672 36168
rect 9864 36159 9916 36168
rect 9864 36125 9873 36159
rect 9873 36125 9907 36159
rect 9907 36125 9916 36159
rect 9864 36116 9916 36125
rect 1952 35980 2004 36032
rect 9864 35980 9916 36032
rect 10048 36023 10100 36032
rect 10048 35989 10057 36023
rect 10057 35989 10091 36023
rect 10091 35989 10100 36023
rect 10048 35980 10100 35989
rect 4213 35878 4265 35930
rect 4277 35878 4329 35930
rect 4341 35878 4393 35930
rect 4405 35878 4457 35930
rect 4469 35878 4521 35930
rect 7477 35878 7529 35930
rect 7541 35878 7593 35930
rect 7605 35878 7657 35930
rect 7669 35878 7721 35930
rect 7733 35878 7785 35930
rect 1676 35683 1728 35692
rect 1676 35649 1685 35683
rect 1685 35649 1719 35683
rect 1719 35649 1728 35683
rect 1676 35640 1728 35649
rect 2412 35776 2464 35828
rect 2504 35776 2556 35828
rect 3332 35776 3384 35828
rect 3608 35776 3660 35828
rect 2596 35640 2648 35692
rect 3332 35640 3384 35692
rect 2044 35572 2096 35624
rect 2320 35547 2372 35556
rect 2320 35513 2329 35547
rect 2329 35513 2363 35547
rect 2363 35513 2372 35547
rect 2320 35504 2372 35513
rect 1492 35479 1544 35488
rect 1492 35445 1501 35479
rect 1501 35445 1535 35479
rect 1535 35445 1544 35479
rect 1492 35436 1544 35445
rect 2582 35334 2634 35386
rect 2646 35334 2698 35386
rect 2710 35334 2762 35386
rect 2774 35334 2826 35386
rect 2838 35334 2890 35386
rect 5845 35334 5897 35386
rect 5909 35334 5961 35386
rect 5973 35334 6025 35386
rect 6037 35334 6089 35386
rect 6101 35334 6153 35386
rect 9109 35334 9161 35386
rect 9173 35334 9225 35386
rect 9237 35334 9289 35386
rect 9301 35334 9353 35386
rect 9365 35334 9417 35386
rect 4620 35096 4672 35148
rect 1952 35028 2004 35080
rect 4804 35028 4856 35080
rect 9864 35071 9916 35080
rect 9864 35037 9873 35071
rect 9873 35037 9907 35071
rect 9907 35037 9916 35071
rect 9864 35028 9916 35037
rect 1584 34935 1636 34944
rect 1584 34901 1593 34935
rect 1593 34901 1627 34935
rect 1627 34901 1636 34935
rect 1584 34892 1636 34901
rect 1676 34892 1728 34944
rect 3700 34892 3752 34944
rect 10048 34935 10100 34944
rect 10048 34901 10057 34935
rect 10057 34901 10091 34935
rect 10091 34901 10100 34935
rect 10048 34892 10100 34901
rect 4213 34790 4265 34842
rect 4277 34790 4329 34842
rect 4341 34790 4393 34842
rect 4405 34790 4457 34842
rect 4469 34790 4521 34842
rect 7477 34790 7529 34842
rect 7541 34790 7593 34842
rect 7605 34790 7657 34842
rect 7669 34790 7721 34842
rect 7733 34790 7785 34842
rect 5080 34688 5132 34740
rect 5448 34620 5500 34672
rect 1860 34552 1912 34604
rect 3056 34595 3108 34604
rect 3056 34561 3065 34595
rect 3065 34561 3099 34595
rect 3099 34561 3108 34595
rect 3056 34552 3108 34561
rect 3240 34484 3292 34536
rect 1492 34348 1544 34400
rect 2582 34246 2634 34298
rect 2646 34246 2698 34298
rect 2710 34246 2762 34298
rect 2774 34246 2826 34298
rect 2838 34246 2890 34298
rect 5845 34246 5897 34298
rect 5909 34246 5961 34298
rect 5973 34246 6025 34298
rect 6037 34246 6089 34298
rect 6101 34246 6153 34298
rect 9109 34246 9161 34298
rect 9173 34246 9225 34298
rect 9237 34246 9289 34298
rect 9301 34246 9353 34298
rect 9365 34246 9417 34298
rect 3056 34187 3108 34196
rect 3056 34153 3065 34187
rect 3065 34153 3099 34187
rect 3099 34153 3108 34187
rect 3056 34144 3108 34153
rect 2044 33940 2096 33992
rect 2320 33983 2372 33992
rect 2320 33949 2329 33983
rect 2329 33949 2363 33983
rect 2363 33949 2372 33983
rect 2320 33940 2372 33949
rect 2412 33940 2464 33992
rect 3056 33940 3108 33992
rect 9864 33983 9916 33992
rect 9864 33949 9873 33983
rect 9873 33949 9907 33983
rect 9907 33949 9916 33983
rect 9864 33940 9916 33949
rect 1584 33847 1636 33856
rect 1584 33813 1593 33847
rect 1593 33813 1627 33847
rect 1627 33813 1636 33847
rect 1584 33804 1636 33813
rect 7288 33872 7340 33924
rect 2872 33804 2924 33856
rect 5632 33804 5684 33856
rect 10048 33847 10100 33856
rect 10048 33813 10057 33847
rect 10057 33813 10091 33847
rect 10091 33813 10100 33847
rect 10048 33804 10100 33813
rect 4213 33702 4265 33754
rect 4277 33702 4329 33754
rect 4341 33702 4393 33754
rect 4405 33702 4457 33754
rect 4469 33702 4521 33754
rect 7477 33702 7529 33754
rect 7541 33702 7593 33754
rect 7605 33702 7657 33754
rect 7669 33702 7721 33754
rect 7733 33702 7785 33754
rect 2872 33600 2924 33652
rect 3148 33643 3200 33652
rect 3148 33609 3157 33643
rect 3157 33609 3191 33643
rect 3191 33609 3200 33643
rect 3148 33600 3200 33609
rect 2412 33532 2464 33584
rect 2044 33464 2096 33516
rect 2320 33507 2372 33516
rect 2320 33473 2329 33507
rect 2329 33473 2363 33507
rect 2363 33473 2372 33507
rect 2320 33464 2372 33473
rect 3148 33507 3200 33516
rect 1860 33396 1912 33448
rect 3148 33473 3157 33507
rect 3157 33473 3191 33507
rect 3191 33473 3200 33507
rect 3148 33464 3200 33473
rect 3424 33507 3476 33516
rect 3424 33473 3433 33507
rect 3433 33473 3467 33507
rect 3467 33473 3476 33507
rect 3424 33464 3476 33473
rect 4252 33464 4304 33516
rect 4528 33507 4580 33516
rect 4528 33473 4537 33507
rect 4537 33473 4571 33507
rect 4571 33473 4580 33507
rect 4528 33464 4580 33473
rect 4896 33328 4948 33380
rect 9864 33260 9916 33312
rect 2582 33158 2634 33210
rect 2646 33158 2698 33210
rect 2710 33158 2762 33210
rect 2774 33158 2826 33210
rect 2838 33158 2890 33210
rect 5845 33158 5897 33210
rect 5909 33158 5961 33210
rect 5973 33158 6025 33210
rect 6037 33158 6089 33210
rect 6101 33158 6153 33210
rect 9109 33158 9161 33210
rect 9173 33158 9225 33210
rect 9237 33158 9289 33210
rect 9301 33158 9353 33210
rect 9365 33158 9417 33210
rect 3240 33056 3292 33108
rect 1584 33031 1636 33040
rect 1584 32997 1593 33031
rect 1593 32997 1627 33031
rect 1627 32997 1636 33031
rect 1584 32988 1636 32997
rect 5356 32988 5408 33040
rect 2504 32920 2556 32972
rect 2320 32852 2372 32904
rect 3240 32895 3292 32904
rect 2780 32784 2832 32836
rect 3240 32861 3249 32895
rect 3249 32861 3283 32895
rect 3283 32861 3292 32895
rect 3240 32852 3292 32861
rect 4252 32852 4304 32904
rect 4528 32895 4580 32904
rect 4528 32861 4537 32895
rect 4537 32861 4571 32895
rect 4571 32861 4580 32895
rect 4528 32852 4580 32861
rect 4896 32784 4948 32836
rect 10048 32759 10100 32768
rect 10048 32725 10057 32759
rect 10057 32725 10091 32759
rect 10091 32725 10100 32759
rect 10048 32716 10100 32725
rect 4213 32614 4265 32666
rect 4277 32614 4329 32666
rect 4341 32614 4393 32666
rect 4405 32614 4457 32666
rect 4469 32614 4521 32666
rect 7477 32614 7529 32666
rect 7541 32614 7593 32666
rect 7605 32614 7657 32666
rect 7669 32614 7721 32666
rect 7733 32614 7785 32666
rect 3516 32512 3568 32564
rect 480 32444 532 32496
rect 3332 32444 3384 32496
rect 1400 32419 1452 32428
rect 1400 32385 1409 32419
rect 1409 32385 1443 32419
rect 1443 32385 1452 32419
rect 1400 32376 1452 32385
rect 2504 32419 2556 32428
rect 2504 32385 2513 32419
rect 2513 32385 2547 32419
rect 2547 32385 2556 32419
rect 4620 32419 4672 32428
rect 2504 32376 2556 32385
rect 4620 32385 4629 32419
rect 4629 32385 4663 32419
rect 4663 32385 4672 32419
rect 4620 32376 4672 32385
rect 2780 32308 2832 32360
rect 3148 32308 3200 32360
rect 4804 32308 4856 32360
rect 2582 32070 2634 32122
rect 2646 32070 2698 32122
rect 2710 32070 2762 32122
rect 2774 32070 2826 32122
rect 2838 32070 2890 32122
rect 5845 32070 5897 32122
rect 5909 32070 5961 32122
rect 5973 32070 6025 32122
rect 6037 32070 6089 32122
rect 6101 32070 6153 32122
rect 9109 32070 9161 32122
rect 9173 32070 9225 32122
rect 9237 32070 9289 32122
rect 9301 32070 9353 32122
rect 9365 32070 9417 32122
rect 1768 31968 1820 32020
rect 2044 31968 2096 32020
rect 3056 31832 3108 31884
rect 2780 31764 2832 31816
rect 4620 31807 4672 31816
rect 1860 31696 1912 31748
rect 4620 31773 4629 31807
rect 4629 31773 4663 31807
rect 4663 31773 4672 31807
rect 4620 31764 4672 31773
rect 10048 31671 10100 31680
rect 10048 31637 10057 31671
rect 10057 31637 10091 31671
rect 10091 31637 10100 31671
rect 10048 31628 10100 31637
rect 4213 31526 4265 31578
rect 4277 31526 4329 31578
rect 4341 31526 4393 31578
rect 4405 31526 4457 31578
rect 4469 31526 4521 31578
rect 7477 31526 7529 31578
rect 7541 31526 7593 31578
rect 7605 31526 7657 31578
rect 7669 31526 7721 31578
rect 7733 31526 7785 31578
rect 2412 31467 2464 31476
rect 2412 31433 2421 31467
rect 2421 31433 2455 31467
rect 2455 31433 2464 31467
rect 2412 31424 2464 31433
rect 3424 31356 3476 31408
rect 2320 31331 2372 31340
rect 2320 31297 2329 31331
rect 2329 31297 2363 31331
rect 2363 31297 2372 31331
rect 2320 31288 2372 31297
rect 2504 31288 2556 31340
rect 4620 31331 4672 31340
rect 4620 31297 4629 31331
rect 4629 31297 4663 31331
rect 4663 31297 4672 31331
rect 4620 31288 4672 31297
rect 3424 31220 3476 31272
rect 9864 31084 9916 31136
rect 2582 30982 2634 31034
rect 2646 30982 2698 31034
rect 2710 30982 2762 31034
rect 2774 30982 2826 31034
rect 2838 30982 2890 31034
rect 5845 30982 5897 31034
rect 5909 30982 5961 31034
rect 5973 30982 6025 31034
rect 6037 30982 6089 31034
rect 6101 30982 6153 31034
rect 9109 30982 9161 31034
rect 9173 30982 9225 31034
rect 9237 30982 9289 31034
rect 9301 30982 9353 31034
rect 9365 30982 9417 31034
rect 1860 30880 1912 30932
rect 2228 30880 2280 30932
rect 3792 30923 3844 30932
rect 3792 30889 3801 30923
rect 3801 30889 3835 30923
rect 3835 30889 3844 30923
rect 3792 30880 3844 30889
rect 2136 30812 2188 30864
rect 1860 30719 1912 30728
rect 1860 30685 1869 30719
rect 1869 30685 1903 30719
rect 1903 30685 1912 30719
rect 1860 30676 1912 30685
rect 2780 30676 2832 30728
rect 3148 30719 3200 30728
rect 3148 30685 3157 30719
rect 3157 30685 3191 30719
rect 3191 30685 3200 30719
rect 3148 30676 3200 30685
rect 3976 30719 4028 30728
rect 3976 30685 3985 30719
rect 3985 30685 4019 30719
rect 4019 30685 4028 30719
rect 3976 30676 4028 30685
rect 4620 30719 4672 30728
rect 4620 30685 4629 30719
rect 4629 30685 4663 30719
rect 4663 30685 4672 30719
rect 4620 30676 4672 30685
rect 9864 30719 9916 30728
rect 9864 30685 9873 30719
rect 9873 30685 9907 30719
rect 9907 30685 9916 30719
rect 9864 30676 9916 30685
rect 4896 30608 4948 30660
rect 9864 30540 9916 30592
rect 10048 30583 10100 30592
rect 10048 30549 10057 30583
rect 10057 30549 10091 30583
rect 10091 30549 10100 30583
rect 10048 30540 10100 30549
rect 4213 30438 4265 30490
rect 4277 30438 4329 30490
rect 4341 30438 4393 30490
rect 4405 30438 4457 30490
rect 4469 30438 4521 30490
rect 7477 30438 7529 30490
rect 7541 30438 7593 30490
rect 7605 30438 7657 30490
rect 7669 30438 7721 30490
rect 7733 30438 7785 30490
rect 2320 30336 2372 30388
rect 2228 30200 2280 30252
rect 2320 30243 2372 30252
rect 2320 30209 2329 30243
rect 2329 30209 2363 30243
rect 2363 30209 2372 30243
rect 2320 30200 2372 30209
rect 2504 30132 2556 30184
rect 2582 29894 2634 29946
rect 2646 29894 2698 29946
rect 2710 29894 2762 29946
rect 2774 29894 2826 29946
rect 2838 29894 2890 29946
rect 5845 29894 5897 29946
rect 5909 29894 5961 29946
rect 5973 29894 6025 29946
rect 6037 29894 6089 29946
rect 6101 29894 6153 29946
rect 9109 29894 9161 29946
rect 9173 29894 9225 29946
rect 9237 29894 9289 29946
rect 9301 29894 9353 29946
rect 9365 29894 9417 29946
rect 1860 29792 1912 29844
rect 3056 29835 3108 29844
rect 3056 29801 3065 29835
rect 3065 29801 3099 29835
rect 3099 29801 3108 29835
rect 3056 29792 3108 29801
rect 4896 29656 4948 29708
rect 2044 29588 2096 29640
rect 3056 29588 3108 29640
rect 3240 29631 3292 29640
rect 3240 29597 3249 29631
rect 3249 29597 3283 29631
rect 3283 29597 3292 29631
rect 3240 29588 3292 29597
rect 9864 29631 9916 29640
rect 9864 29597 9873 29631
rect 9873 29597 9907 29631
rect 9907 29597 9916 29631
rect 9864 29588 9916 29597
rect 10048 29495 10100 29504
rect 10048 29461 10057 29495
rect 10057 29461 10091 29495
rect 10091 29461 10100 29495
rect 10048 29452 10100 29461
rect 4213 29350 4265 29402
rect 4277 29350 4329 29402
rect 4341 29350 4393 29402
rect 4405 29350 4457 29402
rect 4469 29350 4521 29402
rect 7477 29350 7529 29402
rect 7541 29350 7593 29402
rect 7605 29350 7657 29402
rect 7669 29350 7721 29402
rect 7733 29350 7785 29402
rect 2228 29248 2280 29300
rect 3424 29248 3476 29300
rect 6276 29180 6328 29232
rect 1952 29155 2004 29164
rect 1952 29121 1961 29155
rect 1961 29121 1995 29155
rect 1995 29121 2004 29155
rect 1952 29112 2004 29121
rect 1860 29044 1912 29096
rect 3148 29112 3200 29164
rect 3516 29155 3568 29164
rect 3516 29121 3525 29155
rect 3525 29121 3559 29155
rect 3559 29121 3568 29155
rect 3516 29112 3568 29121
rect 3792 29044 3844 29096
rect 2582 28806 2634 28858
rect 2646 28806 2698 28858
rect 2710 28806 2762 28858
rect 2774 28806 2826 28858
rect 2838 28806 2890 28858
rect 5845 28806 5897 28858
rect 5909 28806 5961 28858
rect 5973 28806 6025 28858
rect 6037 28806 6089 28858
rect 6101 28806 6153 28858
rect 9109 28806 9161 28858
rect 9173 28806 9225 28858
rect 9237 28806 9289 28858
rect 9301 28806 9353 28858
rect 9365 28806 9417 28858
rect 3608 28636 3660 28688
rect 572 28568 624 28620
rect 1952 28500 2004 28552
rect 2136 28543 2188 28552
rect 2136 28509 2145 28543
rect 2145 28509 2179 28543
rect 2179 28509 2188 28543
rect 2872 28543 2924 28552
rect 2136 28500 2188 28509
rect 2872 28509 2881 28543
rect 2881 28509 2915 28543
rect 2915 28509 2924 28543
rect 2872 28500 2924 28509
rect 3700 28500 3752 28552
rect 3792 28543 3844 28552
rect 3792 28509 3801 28543
rect 3801 28509 3835 28543
rect 3835 28509 3844 28543
rect 3792 28500 3844 28509
rect 4620 28500 4672 28552
rect 10048 28407 10100 28416
rect 10048 28373 10057 28407
rect 10057 28373 10091 28407
rect 10091 28373 10100 28407
rect 10048 28364 10100 28373
rect 4213 28262 4265 28314
rect 4277 28262 4329 28314
rect 4341 28262 4393 28314
rect 4405 28262 4457 28314
rect 4469 28262 4521 28314
rect 7477 28262 7529 28314
rect 7541 28262 7593 28314
rect 7605 28262 7657 28314
rect 7669 28262 7721 28314
rect 7733 28262 7785 28314
rect 2964 28203 3016 28212
rect 2964 28169 2973 28203
rect 2973 28169 3007 28203
rect 3007 28169 3016 28203
rect 2964 28160 3016 28169
rect 6184 28092 6236 28144
rect 1492 28024 1544 28076
rect 2872 28067 2924 28076
rect 2872 28033 2881 28067
rect 2881 28033 2915 28067
rect 2915 28033 2924 28067
rect 2872 28024 2924 28033
rect 3240 28024 3292 28076
rect 4528 28024 4580 28076
rect 4804 28024 4856 28076
rect 4252 27999 4304 28008
rect 4252 27965 4261 27999
rect 4261 27965 4295 27999
rect 4295 27965 4304 27999
rect 4252 27956 4304 27965
rect 4620 27956 4672 28008
rect 2582 27718 2634 27770
rect 2646 27718 2698 27770
rect 2710 27718 2762 27770
rect 2774 27718 2826 27770
rect 2838 27718 2890 27770
rect 5845 27718 5897 27770
rect 5909 27718 5961 27770
rect 5973 27718 6025 27770
rect 6037 27718 6089 27770
rect 6101 27718 6153 27770
rect 9109 27718 9161 27770
rect 9173 27718 9225 27770
rect 9237 27718 9289 27770
rect 9301 27718 9353 27770
rect 9365 27718 9417 27770
rect 2964 27616 3016 27668
rect 1860 27548 1912 27600
rect 2044 27591 2096 27600
rect 2044 27557 2053 27591
rect 2053 27557 2087 27591
rect 2087 27557 2096 27591
rect 2044 27548 2096 27557
rect 1584 27455 1636 27464
rect 1584 27421 1593 27455
rect 1593 27421 1627 27455
rect 1627 27421 1636 27455
rect 1584 27412 1636 27421
rect 2228 27455 2280 27464
rect 2228 27421 2237 27455
rect 2237 27421 2271 27455
rect 2271 27421 2280 27455
rect 2228 27412 2280 27421
rect 3056 27412 3108 27464
rect 3332 27412 3384 27464
rect 3700 27412 3752 27464
rect 3976 27455 4028 27464
rect 3976 27421 3985 27455
rect 3985 27421 4019 27455
rect 4019 27421 4028 27455
rect 3976 27412 4028 27421
rect 4252 27412 4304 27464
rect 10048 27319 10100 27328
rect 10048 27285 10057 27319
rect 10057 27285 10091 27319
rect 10091 27285 10100 27319
rect 10048 27276 10100 27285
rect 4213 27174 4265 27226
rect 4277 27174 4329 27226
rect 4341 27174 4393 27226
rect 4405 27174 4457 27226
rect 4469 27174 4521 27226
rect 7477 27174 7529 27226
rect 7541 27174 7593 27226
rect 7605 27174 7657 27226
rect 7669 27174 7721 27226
rect 7733 27174 7785 27226
rect 1584 27072 1636 27124
rect 3700 27004 3752 27056
rect 1584 26979 1636 26988
rect 1584 26945 1593 26979
rect 1593 26945 1627 26979
rect 1627 26945 1636 26979
rect 1584 26936 1636 26945
rect 2228 26936 2280 26988
rect 2872 26979 2924 26988
rect 2872 26945 2881 26979
rect 2881 26945 2915 26979
rect 2915 26945 2924 26979
rect 2872 26936 2924 26945
rect 2136 26868 2188 26920
rect 3976 26936 4028 26988
rect 4160 26936 4212 26988
rect 9864 26732 9916 26784
rect 2582 26630 2634 26682
rect 2646 26630 2698 26682
rect 2710 26630 2762 26682
rect 2774 26630 2826 26682
rect 2838 26630 2890 26682
rect 5845 26630 5897 26682
rect 5909 26630 5961 26682
rect 5973 26630 6025 26682
rect 6037 26630 6089 26682
rect 6101 26630 6153 26682
rect 9109 26630 9161 26682
rect 9173 26630 9225 26682
rect 9237 26630 9289 26682
rect 9301 26630 9353 26682
rect 9365 26630 9417 26682
rect 2228 26571 2280 26580
rect 2228 26537 2237 26571
rect 2237 26537 2271 26571
rect 2271 26537 2280 26571
rect 2228 26528 2280 26537
rect 3240 26460 3292 26512
rect 664 26392 716 26444
rect 1860 26324 1912 26376
rect 2044 26367 2096 26376
rect 2044 26333 2053 26367
rect 2053 26333 2087 26367
rect 2087 26333 2096 26367
rect 2044 26324 2096 26333
rect 3792 26367 3844 26376
rect 3792 26333 3801 26367
rect 3801 26333 3835 26367
rect 3835 26333 3844 26367
rect 3792 26324 3844 26333
rect 9956 26460 10008 26512
rect 3240 26256 3292 26308
rect 4160 26256 4212 26308
rect 9864 26367 9916 26376
rect 9864 26333 9873 26367
rect 9873 26333 9907 26367
rect 9907 26333 9916 26367
rect 9864 26324 9916 26333
rect 9772 26256 9824 26308
rect 1492 26188 1544 26240
rect 3792 26188 3844 26240
rect 10048 26231 10100 26240
rect 10048 26197 10057 26231
rect 10057 26197 10091 26231
rect 10091 26197 10100 26231
rect 10048 26188 10100 26197
rect 4213 26086 4265 26138
rect 4277 26086 4329 26138
rect 4341 26086 4393 26138
rect 4405 26086 4457 26138
rect 4469 26086 4521 26138
rect 7477 26086 7529 26138
rect 7541 26086 7593 26138
rect 7605 26086 7657 26138
rect 7669 26086 7721 26138
rect 7733 26086 7785 26138
rect 1492 26027 1544 26036
rect 1492 25993 1501 26027
rect 1501 25993 1535 26027
rect 1535 25993 1544 26027
rect 1492 25984 1544 25993
rect 1584 25984 1636 26036
rect 2044 25848 2096 25900
rect 2228 25891 2280 25900
rect 2228 25857 2237 25891
rect 2237 25857 2271 25891
rect 2271 25857 2280 25891
rect 2228 25848 2280 25857
rect 2582 25542 2634 25594
rect 2646 25542 2698 25594
rect 2710 25542 2762 25594
rect 2774 25542 2826 25594
rect 2838 25542 2890 25594
rect 5845 25542 5897 25594
rect 5909 25542 5961 25594
rect 5973 25542 6025 25594
rect 6037 25542 6089 25594
rect 6101 25542 6153 25594
rect 9109 25542 9161 25594
rect 9173 25542 9225 25594
rect 9237 25542 9289 25594
rect 9301 25542 9353 25594
rect 9365 25542 9417 25594
rect 2044 25483 2096 25492
rect 2044 25449 2053 25483
rect 2053 25449 2087 25483
rect 2087 25449 2096 25483
rect 2044 25440 2096 25449
rect 1860 25372 1912 25424
rect 4068 25304 4120 25356
rect 6368 25304 6420 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 2228 25279 2280 25288
rect 2228 25245 2237 25279
rect 2237 25245 2271 25279
rect 2271 25245 2280 25279
rect 2228 25236 2280 25245
rect 2872 25279 2924 25288
rect 2872 25245 2881 25279
rect 2881 25245 2915 25279
rect 2915 25245 2924 25279
rect 2872 25236 2924 25245
rect 9956 25236 10008 25288
rect 2044 25100 2096 25152
rect 10048 25143 10100 25152
rect 10048 25109 10057 25143
rect 10057 25109 10091 25143
rect 10091 25109 10100 25143
rect 10048 25100 10100 25109
rect 4213 24998 4265 25050
rect 4277 24998 4329 25050
rect 4341 24998 4393 25050
rect 4405 24998 4457 25050
rect 4469 24998 4521 25050
rect 7477 24998 7529 25050
rect 7541 24998 7593 25050
rect 7605 24998 7657 25050
rect 7669 24998 7721 25050
rect 7733 24998 7785 25050
rect 1492 24760 1544 24812
rect 3240 24803 3292 24812
rect 3240 24769 3249 24803
rect 3249 24769 3283 24803
rect 3283 24769 3292 24803
rect 3240 24760 3292 24769
rect 4252 24760 4304 24812
rect 1400 24556 1452 24608
rect 4988 24556 5040 24608
rect 2582 24454 2634 24506
rect 2646 24454 2698 24506
rect 2710 24454 2762 24506
rect 2774 24454 2826 24506
rect 2838 24454 2890 24506
rect 5845 24454 5897 24506
rect 5909 24454 5961 24506
rect 5973 24454 6025 24506
rect 6037 24454 6089 24506
rect 6101 24454 6153 24506
rect 9109 24454 9161 24506
rect 9173 24454 9225 24506
rect 9237 24454 9289 24506
rect 9301 24454 9353 24506
rect 9365 24454 9417 24506
rect 3884 24352 3936 24404
rect 4712 24352 4764 24404
rect 4620 24284 4672 24336
rect 2044 24191 2096 24200
rect 2044 24157 2053 24191
rect 2053 24157 2087 24191
rect 2087 24157 2096 24191
rect 2044 24148 2096 24157
rect 2872 24191 2924 24200
rect 2872 24157 2881 24191
rect 2881 24157 2915 24191
rect 2915 24157 2924 24191
rect 2872 24148 2924 24157
rect 4252 24191 4304 24200
rect 4252 24157 4261 24191
rect 4261 24157 4295 24191
rect 4295 24157 4304 24191
rect 4252 24148 4304 24157
rect 9772 24148 9824 24200
rect 2044 24012 2096 24064
rect 2136 24055 2188 24064
rect 2136 24021 2145 24055
rect 2145 24021 2179 24055
rect 2179 24021 2188 24055
rect 10048 24055 10100 24064
rect 2136 24012 2188 24021
rect 10048 24021 10057 24055
rect 10057 24021 10091 24055
rect 10091 24021 10100 24055
rect 10048 24012 10100 24021
rect 4213 23910 4265 23962
rect 4277 23910 4329 23962
rect 4341 23910 4393 23962
rect 4405 23910 4457 23962
rect 4469 23910 4521 23962
rect 7477 23910 7529 23962
rect 7541 23910 7593 23962
rect 7605 23910 7657 23962
rect 7669 23910 7721 23962
rect 7733 23910 7785 23962
rect 4068 23808 4120 23860
rect 2136 23740 2188 23792
rect 2044 23715 2096 23724
rect 2044 23681 2053 23715
rect 2053 23681 2087 23715
rect 2087 23681 2096 23715
rect 2044 23672 2096 23681
rect 2964 23715 3016 23724
rect 2964 23681 2973 23715
rect 2973 23681 3007 23715
rect 3007 23681 3016 23715
rect 2964 23672 3016 23681
rect 4344 23740 4396 23792
rect 3792 23715 3844 23724
rect 3792 23681 3801 23715
rect 3801 23681 3835 23715
rect 3835 23681 3844 23715
rect 3792 23672 3844 23681
rect 4068 23604 4120 23656
rect 6552 23536 6604 23588
rect 3608 23511 3660 23520
rect 3608 23477 3617 23511
rect 3617 23477 3651 23511
rect 3651 23477 3660 23511
rect 3608 23468 3660 23477
rect 2582 23366 2634 23418
rect 2646 23366 2698 23418
rect 2710 23366 2762 23418
rect 2774 23366 2826 23418
rect 2838 23366 2890 23418
rect 5845 23366 5897 23418
rect 5909 23366 5961 23418
rect 5973 23366 6025 23418
rect 6037 23366 6089 23418
rect 6101 23366 6153 23418
rect 9109 23366 9161 23418
rect 9173 23366 9225 23418
rect 9237 23366 9289 23418
rect 9301 23366 9353 23418
rect 9365 23366 9417 23418
rect 3056 23307 3108 23316
rect 3056 23273 3065 23307
rect 3065 23273 3099 23307
rect 3099 23273 3108 23307
rect 3056 23264 3108 23273
rect 2044 23171 2096 23180
rect 2044 23137 2053 23171
rect 2053 23137 2087 23171
rect 2087 23137 2096 23171
rect 2044 23128 2096 23137
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2964 23128 3016 23180
rect 3148 23060 3200 23112
rect 4068 23103 4120 23112
rect 4068 23069 4077 23103
rect 4077 23069 4111 23103
rect 4111 23069 4120 23103
rect 4068 23060 4120 23069
rect 4620 23128 4672 23180
rect 4344 23060 4396 23112
rect 3424 22992 3476 23044
rect 6644 22992 6696 23044
rect 4712 22924 4764 22976
rect 10048 22967 10100 22976
rect 10048 22933 10057 22967
rect 10057 22933 10091 22967
rect 10091 22933 10100 22967
rect 10048 22924 10100 22933
rect 4213 22822 4265 22874
rect 4277 22822 4329 22874
rect 4341 22822 4393 22874
rect 4405 22822 4457 22874
rect 4469 22822 4521 22874
rect 7477 22822 7529 22874
rect 7541 22822 7593 22874
rect 7605 22822 7657 22874
rect 7669 22822 7721 22874
rect 7733 22822 7785 22874
rect 1768 22720 1820 22772
rect 3884 22720 3936 22772
rect 4712 22720 4764 22772
rect 9864 22720 9916 22772
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 1676 22584 1728 22636
rect 2964 22627 3016 22636
rect 2964 22593 2973 22627
rect 2973 22593 3007 22627
rect 3007 22593 3016 22627
rect 2964 22584 3016 22593
rect 4620 22584 4672 22636
rect 4804 22516 4856 22568
rect 4712 22448 4764 22500
rect 2582 22278 2634 22330
rect 2646 22278 2698 22330
rect 2710 22278 2762 22330
rect 2774 22278 2826 22330
rect 2838 22278 2890 22330
rect 5845 22278 5897 22330
rect 5909 22278 5961 22330
rect 5973 22278 6025 22330
rect 6037 22278 6089 22330
rect 6101 22278 6153 22330
rect 9109 22278 9161 22330
rect 9173 22278 9225 22330
rect 9237 22278 9289 22330
rect 9301 22278 9353 22330
rect 9365 22278 9417 22330
rect 2964 22176 3016 22228
rect 3608 22040 3660 22092
rect 2044 22015 2096 22024
rect 2044 21981 2053 22015
rect 2053 21981 2087 22015
rect 2087 21981 2096 22015
rect 2044 21972 2096 21981
rect 3056 21972 3108 22024
rect 3148 21972 3200 22024
rect 4620 21972 4672 22024
rect 9864 22015 9916 22024
rect 9864 21981 9873 22015
rect 9873 21981 9907 22015
rect 9907 21981 9916 22015
rect 9864 21972 9916 21981
rect 1676 21836 1728 21888
rect 2504 21836 2556 21888
rect 9864 21836 9916 21888
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 4213 21734 4265 21786
rect 4277 21734 4329 21786
rect 4341 21734 4393 21786
rect 4405 21734 4457 21786
rect 4469 21734 4521 21786
rect 7477 21734 7529 21786
rect 7541 21734 7593 21786
rect 7605 21734 7657 21786
rect 7669 21734 7721 21786
rect 7733 21734 7785 21786
rect 1400 21632 1452 21684
rect 1676 21564 1728 21616
rect 1492 21496 1544 21548
rect 1584 21496 1636 21548
rect 2872 21539 2924 21548
rect 2872 21505 2881 21539
rect 2881 21505 2915 21539
rect 2915 21505 2924 21539
rect 2872 21496 2924 21505
rect 3332 21539 3384 21548
rect 3332 21505 3341 21539
rect 3341 21505 3375 21539
rect 3375 21505 3384 21539
rect 3332 21496 3384 21505
rect 4620 21496 4672 21548
rect 4712 21539 4764 21548
rect 4712 21505 4721 21539
rect 4721 21505 4755 21539
rect 4755 21505 4764 21539
rect 4712 21496 4764 21505
rect 1860 21292 1912 21344
rect 2228 21292 2280 21344
rect 3792 21292 3844 21344
rect 4896 21335 4948 21344
rect 4896 21301 4905 21335
rect 4905 21301 4939 21335
rect 4939 21301 4948 21335
rect 4896 21292 4948 21301
rect 2582 21190 2634 21242
rect 2646 21190 2698 21242
rect 2710 21190 2762 21242
rect 2774 21190 2826 21242
rect 2838 21190 2890 21242
rect 5845 21190 5897 21242
rect 5909 21190 5961 21242
rect 5973 21190 6025 21242
rect 6037 21190 6089 21242
rect 6101 21190 6153 21242
rect 9109 21190 9161 21242
rect 9173 21190 9225 21242
rect 9237 21190 9289 21242
rect 9301 21190 9353 21242
rect 9365 21190 9417 21242
rect 4896 21088 4948 21140
rect 9772 21088 9824 21140
rect 4804 20952 4856 21004
rect 1492 20884 1544 20936
rect 1676 20884 1728 20936
rect 3056 20927 3108 20936
rect 3056 20893 3065 20927
rect 3065 20893 3099 20927
rect 3099 20893 3108 20927
rect 3056 20884 3108 20893
rect 4712 20927 4764 20936
rect 4712 20893 4721 20927
rect 4721 20893 4755 20927
rect 4755 20893 4764 20927
rect 4712 20884 4764 20893
rect 9864 20927 9916 20936
rect 9864 20893 9873 20927
rect 9873 20893 9907 20927
rect 9907 20893 9916 20927
rect 9864 20884 9916 20893
rect 1768 20748 1820 20800
rect 2044 20791 2096 20800
rect 2044 20757 2053 20791
rect 2053 20757 2087 20791
rect 2087 20757 2096 20791
rect 2044 20748 2096 20757
rect 3056 20748 3108 20800
rect 10048 20791 10100 20800
rect 10048 20757 10057 20791
rect 10057 20757 10091 20791
rect 10091 20757 10100 20791
rect 10048 20748 10100 20757
rect 4213 20646 4265 20698
rect 4277 20646 4329 20698
rect 4341 20646 4393 20698
rect 4405 20646 4457 20698
rect 4469 20646 4521 20698
rect 7477 20646 7529 20698
rect 7541 20646 7593 20698
rect 7605 20646 7657 20698
rect 7669 20646 7721 20698
rect 7733 20646 7785 20698
rect 4160 20476 4212 20528
rect 1400 20451 1452 20460
rect 1400 20417 1409 20451
rect 1409 20417 1443 20451
rect 1443 20417 1452 20451
rect 1400 20408 1452 20417
rect 2228 20451 2280 20460
rect 2228 20417 2237 20451
rect 2237 20417 2271 20451
rect 2271 20417 2280 20451
rect 2228 20408 2280 20417
rect 2504 20408 2556 20460
rect 3516 20451 3568 20460
rect 3516 20417 3525 20451
rect 3525 20417 3559 20451
rect 3559 20417 3568 20451
rect 3516 20408 3568 20417
rect 2412 20340 2464 20392
rect 7196 20340 7248 20392
rect 4620 20272 4672 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 3332 20247 3384 20256
rect 3332 20213 3341 20247
rect 3341 20213 3375 20247
rect 3375 20213 3384 20247
rect 3332 20204 3384 20213
rect 2582 20102 2634 20154
rect 2646 20102 2698 20154
rect 2710 20102 2762 20154
rect 2774 20102 2826 20154
rect 2838 20102 2890 20154
rect 5845 20102 5897 20154
rect 5909 20102 5961 20154
rect 5973 20102 6025 20154
rect 6037 20102 6089 20154
rect 6101 20102 6153 20154
rect 9109 20102 9161 20154
rect 9173 20102 9225 20154
rect 9237 20102 9289 20154
rect 9301 20102 9353 20154
rect 9365 20102 9417 20154
rect 7104 20000 7156 20052
rect 2964 19932 3016 19984
rect 7012 19932 7064 19984
rect 756 19864 808 19916
rect 2136 19864 2188 19916
rect 3056 19864 3108 19916
rect 3516 19864 3568 19916
rect 5172 19864 5224 19916
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 2504 19839 2556 19848
rect 2504 19805 2513 19839
rect 2513 19805 2547 19839
rect 2547 19805 2556 19839
rect 2504 19796 2556 19805
rect 3148 19796 3200 19848
rect 3792 19839 3844 19848
rect 3792 19805 3801 19839
rect 3801 19805 3835 19839
rect 3835 19805 3844 19839
rect 3792 19796 3844 19805
rect 9772 19796 9824 19848
rect 4988 19728 5040 19780
rect 1860 19660 1912 19712
rect 3056 19660 3108 19712
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 4213 19558 4265 19610
rect 4277 19558 4329 19610
rect 4341 19558 4393 19610
rect 4405 19558 4457 19610
rect 4469 19558 4521 19610
rect 7477 19558 7529 19610
rect 7541 19558 7593 19610
rect 7605 19558 7657 19610
rect 7669 19558 7721 19610
rect 7733 19558 7785 19610
rect 2412 19456 2464 19508
rect 2964 19499 3016 19508
rect 2964 19465 2973 19499
rect 2973 19465 3007 19499
rect 3007 19465 3016 19499
rect 2964 19456 3016 19465
rect 3976 19456 4028 19508
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 2504 19363 2556 19372
rect 2504 19329 2513 19363
rect 2513 19329 2547 19363
rect 2547 19329 2556 19363
rect 4620 19388 4672 19440
rect 2504 19320 2556 19329
rect 4068 19320 4120 19372
rect 4804 19320 4856 19372
rect 2964 19184 3016 19236
rect 3424 19184 3476 19236
rect 2582 19014 2634 19066
rect 2646 19014 2698 19066
rect 2710 19014 2762 19066
rect 2774 19014 2826 19066
rect 2838 19014 2890 19066
rect 5845 19014 5897 19066
rect 5909 19014 5961 19066
rect 5973 19014 6025 19066
rect 6037 19014 6089 19066
rect 6101 19014 6153 19066
rect 9109 19014 9161 19066
rect 9173 19014 9225 19066
rect 9237 19014 9289 19066
rect 9301 19014 9353 19066
rect 9365 19014 9417 19066
rect 3516 18912 3568 18964
rect 2044 18708 2096 18760
rect 2504 18751 2556 18760
rect 2504 18717 2513 18751
rect 2513 18717 2547 18751
rect 2547 18717 2556 18751
rect 2504 18708 2556 18717
rect 3056 18751 3108 18760
rect 3056 18717 3065 18751
rect 3065 18717 3099 18751
rect 3099 18717 3108 18751
rect 3056 18708 3108 18717
rect 3976 18751 4028 18760
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 7840 18640 7892 18692
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 10048 18615 10100 18624
rect 10048 18581 10057 18615
rect 10057 18581 10091 18615
rect 10091 18581 10100 18615
rect 10048 18572 10100 18581
rect 4213 18470 4265 18522
rect 4277 18470 4329 18522
rect 4341 18470 4393 18522
rect 4405 18470 4457 18522
rect 4469 18470 4521 18522
rect 7477 18470 7529 18522
rect 7541 18470 7593 18522
rect 7605 18470 7657 18522
rect 7669 18470 7721 18522
rect 7733 18470 7785 18522
rect 2136 18411 2188 18420
rect 2136 18377 2145 18411
rect 2145 18377 2179 18411
rect 2179 18377 2188 18411
rect 2136 18368 2188 18377
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 1768 18232 1820 18284
rect 3332 18232 3384 18284
rect 3516 18275 3568 18284
rect 3516 18241 3525 18275
rect 3525 18241 3559 18275
rect 3559 18241 3568 18275
rect 3516 18232 3568 18241
rect 4620 18300 4672 18352
rect 4712 18232 4764 18284
rect 3056 18164 3108 18216
rect 848 18096 900 18148
rect 2044 18096 2096 18148
rect 3148 18096 3200 18148
rect 4344 18096 4396 18148
rect 9772 18096 9824 18148
rect 1492 18028 1544 18080
rect 2136 18028 2188 18080
rect 3056 18028 3108 18080
rect 3332 18071 3384 18080
rect 3332 18037 3341 18071
rect 3341 18037 3375 18071
rect 3375 18037 3384 18071
rect 3332 18028 3384 18037
rect 9864 18028 9916 18080
rect 2582 17926 2634 17978
rect 2646 17926 2698 17978
rect 2710 17926 2762 17978
rect 2774 17926 2826 17978
rect 2838 17926 2890 17978
rect 5845 17926 5897 17978
rect 5909 17926 5961 17978
rect 5973 17926 6025 17978
rect 6037 17926 6089 17978
rect 6101 17926 6153 17978
rect 9109 17926 9161 17978
rect 9173 17926 9225 17978
rect 9237 17926 9289 17978
rect 9301 17926 9353 17978
rect 9365 17926 9417 17978
rect 3976 17824 4028 17876
rect 6460 17824 6512 17876
rect 940 17620 992 17672
rect 1584 17620 1636 17672
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 4344 17663 4396 17672
rect 4344 17629 4353 17663
rect 4353 17629 4387 17663
rect 4387 17629 4396 17663
rect 4344 17620 4396 17629
rect 4712 17620 4764 17672
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 9864 17663 9916 17672
rect 9864 17629 9873 17663
rect 9873 17629 9907 17663
rect 9907 17629 9916 17663
rect 9864 17620 9916 17629
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 2228 17484 2280 17536
rect 4988 17484 5040 17536
rect 10048 17527 10100 17536
rect 10048 17493 10057 17527
rect 10057 17493 10091 17527
rect 10091 17493 10100 17527
rect 10048 17484 10100 17493
rect 4213 17382 4265 17434
rect 4277 17382 4329 17434
rect 4341 17382 4393 17434
rect 4405 17382 4457 17434
rect 4469 17382 4521 17434
rect 7477 17382 7529 17434
rect 7541 17382 7593 17434
rect 7605 17382 7657 17434
rect 7669 17382 7721 17434
rect 7733 17382 7785 17434
rect 2044 17280 2096 17332
rect 3700 17280 3752 17332
rect 4988 17280 5040 17332
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 3792 17144 3844 17196
rect 4804 17212 4856 17264
rect 4712 17144 4764 17196
rect 1676 16940 1728 16992
rect 9864 16940 9916 16992
rect 2582 16838 2634 16890
rect 2646 16838 2698 16890
rect 2710 16838 2762 16890
rect 2774 16838 2826 16890
rect 2838 16838 2890 16890
rect 5845 16838 5897 16890
rect 5909 16838 5961 16890
rect 5973 16838 6025 16890
rect 6037 16838 6089 16890
rect 6101 16838 6153 16890
rect 9109 16838 9161 16890
rect 9173 16838 9225 16890
rect 9237 16838 9289 16890
rect 9301 16838 9353 16890
rect 9365 16838 9417 16890
rect 2228 16736 2280 16788
rect 1492 16643 1544 16652
rect 1492 16609 1501 16643
rect 1501 16609 1535 16643
rect 1535 16609 1544 16643
rect 1492 16600 1544 16609
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 3332 16532 3384 16584
rect 9772 16532 9824 16584
rect 2136 16439 2188 16448
rect 2136 16405 2145 16439
rect 2145 16405 2179 16439
rect 2179 16405 2188 16439
rect 2136 16396 2188 16405
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 4213 16294 4265 16346
rect 4277 16294 4329 16346
rect 4341 16294 4393 16346
rect 4405 16294 4457 16346
rect 4469 16294 4521 16346
rect 7477 16294 7529 16346
rect 7541 16294 7593 16346
rect 7605 16294 7657 16346
rect 7669 16294 7721 16346
rect 7733 16294 7785 16346
rect 1492 16056 1544 16108
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 1952 15920 2004 15972
rect 1860 15852 1912 15904
rect 2582 15750 2634 15802
rect 2646 15750 2698 15802
rect 2710 15750 2762 15802
rect 2774 15750 2826 15802
rect 2838 15750 2890 15802
rect 5845 15750 5897 15802
rect 5909 15750 5961 15802
rect 5973 15750 6025 15802
rect 6037 15750 6089 15802
rect 6101 15750 6153 15802
rect 9109 15750 9161 15802
rect 9173 15750 9225 15802
rect 9237 15750 9289 15802
rect 9301 15750 9353 15802
rect 9365 15750 9417 15802
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 2044 15351 2096 15360
rect 2044 15317 2053 15351
rect 2053 15317 2087 15351
rect 2087 15317 2096 15351
rect 2044 15308 2096 15317
rect 10048 15351 10100 15360
rect 10048 15317 10057 15351
rect 10057 15317 10091 15351
rect 10091 15317 10100 15351
rect 10048 15308 10100 15317
rect 4213 15206 4265 15258
rect 4277 15206 4329 15258
rect 4341 15206 4393 15258
rect 4405 15206 4457 15258
rect 4469 15206 4521 15258
rect 7477 15206 7529 15258
rect 7541 15206 7593 15258
rect 7605 15206 7657 15258
rect 7669 15206 7721 15258
rect 7733 15206 7785 15258
rect 2044 15036 2096 15088
rect 1676 14968 1728 15020
rect 1768 14807 1820 14816
rect 1768 14773 1777 14807
rect 1777 14773 1811 14807
rect 1811 14773 1820 14807
rect 1768 14764 1820 14773
rect 2582 14662 2634 14714
rect 2646 14662 2698 14714
rect 2710 14662 2762 14714
rect 2774 14662 2826 14714
rect 2838 14662 2890 14714
rect 5845 14662 5897 14714
rect 5909 14662 5961 14714
rect 5973 14662 6025 14714
rect 6037 14662 6089 14714
rect 6101 14662 6153 14714
rect 9109 14662 9161 14714
rect 9173 14662 9225 14714
rect 9237 14662 9289 14714
rect 9301 14662 9353 14714
rect 9365 14662 9417 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 2412 14492 2464 14544
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 2136 14356 2188 14408
rect 2320 14399 2372 14408
rect 2320 14365 2329 14399
rect 2329 14365 2363 14399
rect 2363 14365 2372 14399
rect 2320 14356 2372 14365
rect 1952 14288 2004 14340
rect 2136 14220 2188 14272
rect 2504 14263 2556 14272
rect 2504 14229 2513 14263
rect 2513 14229 2547 14263
rect 2547 14229 2556 14263
rect 2504 14220 2556 14229
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 4213 14118 4265 14170
rect 4277 14118 4329 14170
rect 4341 14118 4393 14170
rect 4405 14118 4457 14170
rect 4469 14118 4521 14170
rect 7477 14118 7529 14170
rect 7541 14118 7593 14170
rect 7605 14118 7657 14170
rect 7669 14118 7721 14170
rect 7733 14118 7785 14170
rect 1676 14016 1728 14068
rect 1952 14016 2004 14068
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 2582 13574 2634 13626
rect 2646 13574 2698 13626
rect 2710 13574 2762 13626
rect 2774 13574 2826 13626
rect 2838 13574 2890 13626
rect 5845 13574 5897 13626
rect 5909 13574 5961 13626
rect 5973 13574 6025 13626
rect 6037 13574 6089 13626
rect 6101 13574 6153 13626
rect 9109 13574 9161 13626
rect 9173 13574 9225 13626
rect 9237 13574 9289 13626
rect 9301 13574 9353 13626
rect 9365 13574 9417 13626
rect 1492 13268 1544 13320
rect 1768 13132 1820 13184
rect 4213 13030 4265 13082
rect 4277 13030 4329 13082
rect 4341 13030 4393 13082
rect 4405 13030 4457 13082
rect 4469 13030 4521 13082
rect 7477 13030 7529 13082
rect 7541 13030 7593 13082
rect 7605 13030 7657 13082
rect 7669 13030 7721 13082
rect 7733 13030 7785 13082
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 2228 12835 2280 12844
rect 2228 12801 2237 12835
rect 2237 12801 2271 12835
rect 2271 12801 2280 12835
rect 2228 12792 2280 12801
rect 10048 12699 10100 12708
rect 10048 12665 10057 12699
rect 10057 12665 10091 12699
rect 10091 12665 10100 12699
rect 10048 12656 10100 12665
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 2582 12486 2634 12538
rect 2646 12486 2698 12538
rect 2710 12486 2762 12538
rect 2774 12486 2826 12538
rect 2838 12486 2890 12538
rect 5845 12486 5897 12538
rect 5909 12486 5961 12538
rect 5973 12486 6025 12538
rect 6037 12486 6089 12538
rect 6101 12486 6153 12538
rect 9109 12486 9161 12538
rect 9173 12486 9225 12538
rect 9237 12486 9289 12538
rect 9301 12486 9353 12538
rect 9365 12486 9417 12538
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 1860 12180 1912 12232
rect 1676 12112 1728 12164
rect 1584 12044 1636 12096
rect 1860 12044 1912 12096
rect 4213 11942 4265 11994
rect 4277 11942 4329 11994
rect 4341 11942 4393 11994
rect 4405 11942 4457 11994
rect 4469 11942 4521 11994
rect 7477 11942 7529 11994
rect 7541 11942 7593 11994
rect 7605 11942 7657 11994
rect 7669 11942 7721 11994
rect 7733 11942 7785 11994
rect 2412 11772 2464 11824
rect 1860 11704 1912 11756
rect 2136 11704 2188 11756
rect 3424 11704 3476 11756
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 2044 11636 2096 11688
rect 1952 11568 2004 11620
rect 1768 11500 1820 11552
rect 2044 11500 2096 11552
rect 2504 11636 2556 11688
rect 10048 11611 10100 11620
rect 10048 11577 10057 11611
rect 10057 11577 10091 11611
rect 10091 11577 10100 11611
rect 10048 11568 10100 11577
rect 2320 11500 2372 11552
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 2582 11398 2634 11450
rect 2646 11398 2698 11450
rect 2710 11398 2762 11450
rect 2774 11398 2826 11450
rect 2838 11398 2890 11450
rect 5845 11398 5897 11450
rect 5909 11398 5961 11450
rect 5973 11398 6025 11450
rect 6037 11398 6089 11450
rect 6101 11398 6153 11450
rect 9109 11398 9161 11450
rect 9173 11398 9225 11450
rect 9237 11398 9289 11450
rect 9301 11398 9353 11450
rect 9365 11398 9417 11450
rect 1676 11296 1728 11348
rect 2504 11296 2556 11348
rect 2964 11160 3016 11212
rect 3884 11160 3936 11212
rect 5264 11160 5316 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 3056 11092 3108 11144
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 4620 11092 4672 11144
rect 112 11024 164 11076
rect 2964 11024 3016 11076
rect 9864 11024 9916 11076
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 4213 10854 4265 10906
rect 4277 10854 4329 10906
rect 4341 10854 4393 10906
rect 4405 10854 4457 10906
rect 4469 10854 4521 10906
rect 7477 10854 7529 10906
rect 7541 10854 7593 10906
rect 7605 10854 7657 10906
rect 7669 10854 7721 10906
rect 7733 10854 7785 10906
rect 3240 10752 3292 10804
rect 2136 10684 2188 10736
rect 1860 10616 1912 10668
rect 2320 10616 2372 10668
rect 4896 10616 4948 10668
rect 9864 10659 9916 10668
rect 9864 10625 9873 10659
rect 9873 10625 9907 10659
rect 9907 10625 9916 10659
rect 9864 10616 9916 10625
rect 4620 10591 4672 10600
rect 4620 10557 4629 10591
rect 4629 10557 4663 10591
rect 4663 10557 4672 10591
rect 4620 10548 4672 10557
rect 10048 10523 10100 10532
rect 10048 10489 10057 10523
rect 10057 10489 10091 10523
rect 10091 10489 10100 10523
rect 10048 10480 10100 10489
rect 2582 10310 2634 10362
rect 2646 10310 2698 10362
rect 2710 10310 2762 10362
rect 2774 10310 2826 10362
rect 2838 10310 2890 10362
rect 5845 10310 5897 10362
rect 5909 10310 5961 10362
rect 5973 10310 6025 10362
rect 6037 10310 6089 10362
rect 6101 10310 6153 10362
rect 9109 10310 9161 10362
rect 9173 10310 9225 10362
rect 9237 10310 9289 10362
rect 9301 10310 9353 10362
rect 9365 10310 9417 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 2228 10208 2280 10260
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 2044 10004 2096 10056
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 4620 10004 4672 10056
rect 1032 9936 1084 9988
rect 2228 9936 2280 9988
rect 9864 9868 9916 9920
rect 4213 9766 4265 9818
rect 4277 9766 4329 9818
rect 4341 9766 4393 9818
rect 4405 9766 4457 9818
rect 4469 9766 4521 9818
rect 7477 9766 7529 9818
rect 7541 9766 7593 9818
rect 7605 9766 7657 9818
rect 7669 9766 7721 9818
rect 7733 9766 7785 9818
rect 9864 9664 9916 9716
rect 3700 9528 3752 9580
rect 4620 9528 4672 9580
rect 4896 9528 4948 9580
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 10048 9435 10100 9444
rect 10048 9401 10057 9435
rect 10057 9401 10091 9435
rect 10091 9401 10100 9435
rect 10048 9392 10100 9401
rect 9864 9324 9916 9376
rect 2582 9222 2634 9274
rect 2646 9222 2698 9274
rect 2710 9222 2762 9274
rect 2774 9222 2826 9274
rect 2838 9222 2890 9274
rect 5845 9222 5897 9274
rect 5909 9222 5961 9274
rect 5973 9222 6025 9274
rect 6037 9222 6089 9274
rect 6101 9222 6153 9274
rect 9109 9222 9161 9274
rect 9173 9222 9225 9274
rect 9237 9222 9289 9274
rect 9301 9222 9353 9274
rect 9365 9222 9417 9274
rect 4213 8678 4265 8730
rect 4277 8678 4329 8730
rect 4341 8678 4393 8730
rect 4405 8678 4457 8730
rect 4469 8678 4521 8730
rect 7477 8678 7529 8730
rect 7541 8678 7593 8730
rect 7605 8678 7657 8730
rect 7669 8678 7721 8730
rect 7733 8678 7785 8730
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10048 8347 10100 8356
rect 10048 8313 10057 8347
rect 10057 8313 10091 8347
rect 10091 8313 10100 8347
rect 10048 8304 10100 8313
rect 2582 8134 2634 8186
rect 2646 8134 2698 8186
rect 2710 8134 2762 8186
rect 2774 8134 2826 8186
rect 2838 8134 2890 8186
rect 5845 8134 5897 8186
rect 5909 8134 5961 8186
rect 5973 8134 6025 8186
rect 6037 8134 6089 8186
rect 6101 8134 6153 8186
rect 9109 8134 9161 8186
rect 9173 8134 9225 8186
rect 9237 8134 9289 8186
rect 9301 8134 9353 8186
rect 9365 8134 9417 8186
rect 3884 7871 3936 7880
rect 3884 7837 3893 7871
rect 3893 7837 3927 7871
rect 3927 7837 3936 7871
rect 3884 7828 3936 7837
rect 4620 7828 4672 7880
rect 9864 7692 9916 7744
rect 4213 7590 4265 7642
rect 4277 7590 4329 7642
rect 4341 7590 4393 7642
rect 4405 7590 4457 7642
rect 4469 7590 4521 7642
rect 7477 7590 7529 7642
rect 7541 7590 7593 7642
rect 7605 7590 7657 7642
rect 7669 7590 7721 7642
rect 7733 7590 7785 7642
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 10048 7259 10100 7268
rect 10048 7225 10057 7259
rect 10057 7225 10091 7259
rect 10091 7225 10100 7259
rect 10048 7216 10100 7225
rect 2582 7046 2634 7098
rect 2646 7046 2698 7098
rect 2710 7046 2762 7098
rect 2774 7046 2826 7098
rect 2838 7046 2890 7098
rect 5845 7046 5897 7098
rect 5909 7046 5961 7098
rect 5973 7046 6025 7098
rect 6037 7046 6089 7098
rect 6101 7046 6153 7098
rect 9109 7046 9161 7098
rect 9173 7046 9225 7098
rect 9237 7046 9289 7098
rect 9301 7046 9353 7098
rect 9365 7046 9417 7098
rect 2964 6740 3016 6792
rect 5080 6740 5132 6792
rect 9864 6604 9916 6656
rect 4213 6502 4265 6554
rect 4277 6502 4329 6554
rect 4341 6502 4393 6554
rect 4405 6502 4457 6554
rect 4469 6502 4521 6554
rect 7477 6502 7529 6554
rect 7541 6502 7593 6554
rect 7605 6502 7657 6554
rect 7669 6502 7721 6554
rect 7733 6502 7785 6554
rect 3884 6400 3936 6452
rect 2228 6375 2280 6384
rect 2228 6341 2237 6375
rect 2237 6341 2271 6375
rect 2271 6341 2280 6375
rect 2228 6332 2280 6341
rect 1676 6264 1728 6316
rect 3148 6264 3200 6316
rect 5080 6264 5132 6316
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 3884 6128 3936 6180
rect 6828 6128 6880 6180
rect 9772 6060 9824 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 2582 5958 2634 6010
rect 2646 5958 2698 6010
rect 2710 5958 2762 6010
rect 2774 5958 2826 6010
rect 2838 5958 2890 6010
rect 5845 5958 5897 6010
rect 5909 5958 5961 6010
rect 5973 5958 6025 6010
rect 6037 5958 6089 6010
rect 6101 5958 6153 6010
rect 9109 5958 9161 6010
rect 9173 5958 9225 6010
rect 9237 5958 9289 6010
rect 9301 5958 9353 6010
rect 9365 5958 9417 6010
rect 1216 5856 1268 5908
rect 3884 5856 3936 5908
rect 1492 5652 1544 5704
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 3056 5652 3108 5704
rect 5080 5652 5132 5704
rect 5356 5652 5408 5704
rect 1124 5516 1176 5568
rect 9864 5516 9916 5568
rect 4213 5414 4265 5466
rect 4277 5414 4329 5466
rect 4341 5414 4393 5466
rect 4405 5414 4457 5466
rect 4469 5414 4521 5466
rect 7477 5414 7529 5466
rect 7541 5414 7593 5466
rect 7605 5414 7657 5466
rect 7669 5414 7721 5466
rect 7733 5414 7785 5466
rect 1308 5312 1360 5364
rect 2964 5312 3016 5364
rect 1584 5176 1636 5228
rect 2964 5176 3016 5228
rect 5080 5176 5132 5228
rect 9772 5176 9824 5228
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 2582 4870 2634 4922
rect 2646 4870 2698 4922
rect 2710 4870 2762 4922
rect 2774 4870 2826 4922
rect 2838 4870 2890 4922
rect 5845 4870 5897 4922
rect 5909 4870 5961 4922
rect 5973 4870 6025 4922
rect 6037 4870 6089 4922
rect 6101 4870 6153 4922
rect 9109 4870 9161 4922
rect 9173 4870 9225 4922
rect 9237 4870 9289 4922
rect 9301 4870 9353 4922
rect 9365 4870 9417 4922
rect 3148 4768 3200 4820
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 4213 4326 4265 4378
rect 4277 4326 4329 4378
rect 4341 4326 4393 4378
rect 4405 4326 4457 4378
rect 4469 4326 4521 4378
rect 7477 4326 7529 4378
rect 7541 4326 7593 4378
rect 7605 4326 7657 4378
rect 7669 4326 7721 4378
rect 7733 4326 7785 4378
rect 4804 4156 4856 4208
rect 1216 4088 1268 4140
rect 2964 3952 3016 4004
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 2582 3782 2634 3834
rect 2646 3782 2698 3834
rect 2710 3782 2762 3834
rect 2774 3782 2826 3834
rect 2838 3782 2890 3834
rect 5845 3782 5897 3834
rect 5909 3782 5961 3834
rect 5973 3782 6025 3834
rect 6037 3782 6089 3834
rect 6101 3782 6153 3834
rect 9109 3782 9161 3834
rect 9173 3782 9225 3834
rect 9237 3782 9289 3834
rect 9301 3782 9353 3834
rect 9365 3782 9417 3834
rect 1676 3680 1728 3732
rect 1308 3476 1360 3528
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 10048 3383 10100 3392
rect 10048 3349 10057 3383
rect 10057 3349 10091 3383
rect 10091 3349 10100 3383
rect 10048 3340 10100 3349
rect 4213 3238 4265 3290
rect 4277 3238 4329 3290
rect 4341 3238 4393 3290
rect 4405 3238 4457 3290
rect 4469 3238 4521 3290
rect 7477 3238 7529 3290
rect 7541 3238 7593 3290
rect 7605 3238 7657 3290
rect 7669 3238 7721 3290
rect 7733 3238 7785 3290
rect 1584 3179 1636 3188
rect 1584 3145 1593 3179
rect 1593 3145 1627 3179
rect 1627 3145 1636 3179
rect 1584 3136 1636 3145
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 2582 2694 2634 2746
rect 2646 2694 2698 2746
rect 2710 2694 2762 2746
rect 2774 2694 2826 2746
rect 2838 2694 2890 2746
rect 5845 2694 5897 2746
rect 5909 2694 5961 2746
rect 5973 2694 6025 2746
rect 6037 2694 6089 2746
rect 6101 2694 6153 2746
rect 9109 2694 9161 2746
rect 9173 2694 9225 2746
rect 9237 2694 9289 2746
rect 9301 2694 9353 2746
rect 9365 2694 9417 2746
rect 1492 2592 1544 2644
rect 2136 2592 2188 2644
rect 2964 2592 3016 2644
rect 1308 2388 1360 2440
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 2780 2388 2832 2440
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 4213 2150 4265 2202
rect 4277 2150 4329 2202
rect 4341 2150 4393 2202
rect 4405 2150 4457 2202
rect 4469 2150 4521 2202
rect 7477 2150 7529 2202
rect 7541 2150 7593 2202
rect 7605 2150 7657 2202
rect 7669 2150 7721 2202
rect 7733 2150 7785 2202
rect 10968 663 11020 672
rect 10968 629 10977 663
rect 10977 629 11011 663
rect 11011 629 11020 663
rect 10968 620 11020 629
<< metal2 >>
rect 3146 79656 3202 79665
rect 3146 79591 3202 79600
rect 3054 79248 3110 79257
rect 3054 79183 3110 79192
rect 2962 78296 3018 78305
rect 2962 78231 3018 78240
rect 2582 77820 2890 77840
rect 2582 77818 2588 77820
rect 2644 77818 2668 77820
rect 2724 77818 2748 77820
rect 2804 77818 2828 77820
rect 2884 77818 2890 77820
rect 2644 77766 2646 77818
rect 2826 77766 2828 77818
rect 2582 77764 2588 77766
rect 2644 77764 2668 77766
rect 2724 77764 2748 77766
rect 2804 77764 2828 77766
rect 2884 77764 2890 77766
rect 2582 77744 2890 77764
rect 2870 77616 2926 77625
rect 2870 77551 2926 77560
rect 2884 77518 2912 77551
rect 1492 77512 1544 77518
rect 2044 77512 2096 77518
rect 1492 77454 1544 77460
rect 2042 77480 2044 77489
rect 2872 77512 2924 77518
rect 2096 77480 2098 77489
rect 1400 77036 1452 77042
rect 1400 76978 1452 76984
rect 1308 76424 1360 76430
rect 1308 76366 1360 76372
rect 1124 75472 1176 75478
rect 1124 75414 1176 75420
rect 940 75268 992 75274
rect 940 75210 992 75216
rect 952 74866 980 75210
rect 940 74860 992 74866
rect 940 74802 992 74808
rect 388 71120 440 71126
rect 388 71062 440 71068
rect 20 64592 72 64598
rect 20 64534 72 64540
rect 32 42838 60 64534
rect 296 61804 348 61810
rect 296 61746 348 61752
rect 308 55162 336 61746
rect 124 55134 336 55162
rect 124 46170 152 55134
rect 296 52624 348 52630
rect 296 52566 348 52572
rect 204 49700 256 49706
rect 204 49642 256 49648
rect 216 46782 244 49642
rect 204 46776 256 46782
rect 204 46718 256 46724
rect 204 46640 256 46646
rect 204 46582 256 46588
rect 112 46164 164 46170
rect 112 46106 164 46112
rect 112 44464 164 44470
rect 112 44406 164 44412
rect 20 42832 72 42838
rect 20 42774 72 42780
rect 20 42696 72 42702
rect 20 42638 72 42644
rect 32 35894 60 42638
rect 124 40730 152 44406
rect 216 41414 244 46582
rect 308 46238 336 52566
rect 296 46232 348 46238
rect 296 46174 348 46180
rect 296 46096 348 46102
rect 296 46038 348 46044
rect 308 42430 336 46038
rect 400 45626 428 71062
rect 848 69964 900 69970
rect 848 69906 900 69912
rect 664 66496 716 66502
rect 664 66438 716 66444
rect 480 60716 532 60722
rect 480 60658 532 60664
rect 388 45620 440 45626
rect 388 45562 440 45568
rect 296 42424 348 42430
rect 296 42366 348 42372
rect 216 41386 336 41414
rect 112 40724 164 40730
rect 112 40666 164 40672
rect 308 40662 336 41386
rect 296 40656 348 40662
rect 296 40598 348 40604
rect 32 35866 152 35894
rect 124 11082 152 35866
rect 492 32502 520 60658
rect 572 59628 624 59634
rect 572 59570 624 59576
rect 480 32496 532 32502
rect 480 32438 532 32444
rect 584 28626 612 59570
rect 676 56710 704 66438
rect 756 65476 808 65482
rect 756 65418 808 65424
rect 768 56914 796 65418
rect 756 56908 808 56914
rect 756 56850 808 56856
rect 664 56704 716 56710
rect 664 56646 716 56652
rect 664 54664 716 54670
rect 664 54606 716 54612
rect 676 47802 704 54606
rect 860 52494 888 69906
rect 952 64870 980 74802
rect 1032 72208 1084 72214
rect 1032 72150 1084 72156
rect 940 64864 992 64870
rect 940 64806 992 64812
rect 940 63980 992 63986
rect 940 63922 992 63928
rect 848 52488 900 52494
rect 848 52430 900 52436
rect 756 48204 808 48210
rect 756 48146 808 48152
rect 664 47796 716 47802
rect 664 47738 716 47744
rect 664 46232 716 46238
rect 664 46174 716 46180
rect 572 28620 624 28626
rect 572 28562 624 28568
rect 676 26450 704 46174
rect 768 42702 796 48146
rect 848 47524 900 47530
rect 848 47466 900 47472
rect 860 44470 888 47466
rect 848 44464 900 44470
rect 848 44406 900 44412
rect 952 42770 980 63922
rect 1044 47122 1072 72150
rect 1136 49298 1164 75414
rect 1320 75177 1348 76366
rect 1412 76129 1440 76978
rect 1504 76537 1532 77454
rect 2872 77454 2924 77460
rect 2042 77415 2098 77424
rect 1584 77376 1636 77382
rect 1584 77318 1636 77324
rect 2136 77376 2188 77382
rect 2136 77318 2188 77324
rect 2412 77376 2464 77382
rect 2412 77318 2464 77324
rect 2872 77376 2924 77382
rect 2872 77318 2924 77324
rect 1490 76528 1546 76537
rect 1490 76463 1546 76472
rect 1398 76120 1454 76129
rect 1398 76055 1454 76064
rect 1400 75948 1452 75954
rect 1400 75890 1452 75896
rect 1492 75948 1544 75954
rect 1492 75890 1544 75896
rect 1306 75168 1362 75177
rect 1306 75103 1362 75112
rect 1412 74361 1440 75890
rect 1398 74352 1454 74361
rect 1398 74287 1454 74296
rect 1308 74248 1360 74254
rect 1308 74190 1360 74196
rect 1320 73409 1348 74190
rect 1400 73772 1452 73778
rect 1400 73714 1452 73720
rect 1306 73400 1362 73409
rect 1306 73335 1362 73344
rect 1308 73160 1360 73166
rect 1308 73102 1360 73108
rect 1216 72684 1268 72690
rect 1216 72626 1268 72632
rect 1228 71641 1256 72626
rect 1320 72049 1348 73102
rect 1412 73001 1440 73714
rect 1398 72992 1454 73001
rect 1398 72927 1454 72936
rect 1504 72078 1532 75890
rect 1400 72072 1452 72078
rect 1306 72040 1362 72049
rect 1400 72014 1452 72020
rect 1492 72072 1544 72078
rect 1492 72014 1544 72020
rect 1306 71975 1362 71984
rect 1214 71632 1270 71641
rect 1214 71567 1270 71576
rect 1308 71596 1360 71602
rect 1308 71538 1360 71544
rect 1216 70440 1268 70446
rect 1216 70382 1268 70388
rect 1228 69329 1256 70382
rect 1320 70281 1348 71538
rect 1412 71097 1440 72014
rect 1492 71936 1544 71942
rect 1492 71878 1544 71884
rect 1398 71088 1454 71097
rect 1398 71023 1454 71032
rect 1400 70984 1452 70990
rect 1400 70926 1452 70932
rect 1412 70582 1440 70926
rect 1400 70576 1452 70582
rect 1400 70518 1452 70524
rect 1306 70272 1362 70281
rect 1306 70207 1362 70216
rect 1412 70038 1440 70518
rect 1400 70032 1452 70038
rect 1400 69974 1452 69980
rect 1400 69896 1452 69902
rect 1400 69838 1452 69844
rect 1308 69352 1360 69358
rect 1214 69320 1270 69329
rect 1308 69294 1360 69300
rect 1214 69255 1270 69264
rect 1320 68513 1348 69294
rect 1412 68921 1440 69838
rect 1398 68912 1454 68921
rect 1398 68847 1454 68856
rect 1400 68808 1452 68814
rect 1400 68750 1452 68756
rect 1306 68504 1362 68513
rect 1306 68439 1362 68448
rect 1412 67969 1440 68750
rect 1504 68270 1532 71878
rect 1596 71670 1624 77318
rect 2044 77036 2096 77042
rect 2044 76978 2096 76984
rect 2056 76945 2084 76978
rect 2042 76936 2098 76945
rect 2042 76871 2098 76880
rect 1676 76832 1728 76838
rect 1676 76774 1728 76780
rect 1688 75954 1716 76774
rect 2044 76288 2096 76294
rect 2044 76230 2096 76236
rect 1860 76084 1912 76090
rect 1860 76026 1912 76032
rect 1952 76084 2004 76090
rect 1952 76026 2004 76032
rect 1676 75948 1728 75954
rect 1676 75890 1728 75896
rect 1676 74112 1728 74118
rect 1676 74054 1728 74060
rect 1584 71664 1636 71670
rect 1584 71606 1636 71612
rect 1584 71392 1636 71398
rect 1584 71334 1636 71340
rect 1596 70394 1624 71334
rect 1688 70553 1716 74054
rect 1872 72826 1900 76026
rect 1860 72820 1912 72826
rect 1860 72762 1912 72768
rect 1768 72480 1820 72486
rect 1768 72422 1820 72428
rect 1860 72480 1912 72486
rect 1860 72422 1912 72428
rect 1674 70544 1730 70553
rect 1674 70479 1730 70488
rect 1596 70366 1716 70394
rect 1584 70032 1636 70038
rect 1584 69974 1636 69980
rect 1596 68950 1624 69974
rect 1584 68944 1636 68950
rect 1584 68886 1636 68892
rect 1584 68808 1636 68814
rect 1584 68750 1636 68756
rect 1492 68264 1544 68270
rect 1492 68206 1544 68212
rect 1492 68128 1544 68134
rect 1492 68070 1544 68076
rect 1398 67960 1454 67969
rect 1504 67930 1532 68070
rect 1398 67895 1454 67904
rect 1492 67924 1544 67930
rect 1492 67866 1544 67872
rect 1490 67824 1546 67833
rect 1490 67759 1546 67768
rect 1398 67552 1454 67561
rect 1398 67487 1454 67496
rect 1412 67250 1440 67487
rect 1400 67244 1452 67250
rect 1400 67186 1452 67192
rect 1400 66564 1452 66570
rect 1400 66506 1452 66512
rect 1412 66201 1440 66506
rect 1398 66192 1454 66201
rect 1398 66127 1454 66136
rect 1504 66042 1532 67759
rect 1412 66014 1532 66042
rect 1412 64054 1440 66014
rect 1492 64932 1544 64938
rect 1492 64874 1544 64880
rect 1400 64048 1452 64054
rect 1400 63990 1452 63996
rect 1400 63776 1452 63782
rect 1400 63718 1452 63724
rect 1412 62665 1440 63718
rect 1504 63481 1532 64874
rect 1490 63472 1546 63481
rect 1490 63407 1546 63416
rect 1492 63232 1544 63238
rect 1492 63174 1544 63180
rect 1398 62656 1454 62665
rect 1398 62591 1454 62600
rect 1400 62144 1452 62150
rect 1504 62121 1532 63174
rect 1400 62086 1452 62092
rect 1490 62112 1546 62121
rect 1412 61305 1440 62086
rect 1490 62047 1546 62056
rect 1492 61600 1544 61606
rect 1492 61542 1544 61548
rect 1398 61296 1454 61305
rect 1398 61231 1454 61240
rect 1400 61056 1452 61062
rect 1400 60998 1452 61004
rect 1412 60353 1440 60998
rect 1504 60761 1532 61542
rect 1490 60752 1546 60761
rect 1490 60687 1546 60696
rect 1492 60512 1544 60518
rect 1492 60454 1544 60460
rect 1398 60344 1454 60353
rect 1398 60279 1454 60288
rect 1400 59968 1452 59974
rect 1504 59945 1532 60454
rect 1400 59910 1452 59916
rect 1490 59936 1546 59945
rect 1412 58993 1440 59910
rect 1490 59871 1546 59880
rect 1492 59424 1544 59430
rect 1492 59366 1544 59372
rect 1398 58984 1454 58993
rect 1398 58919 1454 58928
rect 1400 58880 1452 58886
rect 1400 58822 1452 58828
rect 1412 58546 1440 58822
rect 1400 58540 1452 58546
rect 1400 58482 1452 58488
rect 1412 58018 1440 58482
rect 1504 58177 1532 59366
rect 1596 58562 1624 68750
rect 1688 68218 1716 70366
rect 1780 68678 1808 72422
rect 1768 68672 1820 68678
rect 1768 68614 1820 68620
rect 1872 68474 1900 72422
rect 1964 70922 1992 76026
rect 2056 75342 2084 76230
rect 2044 75336 2096 75342
rect 2044 75278 2096 75284
rect 2148 73098 2176 77318
rect 2320 76832 2372 76838
rect 2320 76774 2372 76780
rect 2228 75948 2280 75954
rect 2228 75890 2280 75896
rect 2240 75585 2268 75890
rect 2226 75576 2282 75585
rect 2226 75511 2282 75520
rect 2332 75426 2360 76774
rect 2240 75398 2360 75426
rect 2136 73092 2188 73098
rect 2136 73034 2188 73040
rect 2136 72820 2188 72826
rect 2136 72762 2188 72768
rect 2044 72684 2096 72690
rect 2044 72626 2096 72632
rect 2056 72457 2084 72626
rect 2042 72448 2098 72457
rect 2042 72383 2098 72392
rect 2044 72072 2096 72078
rect 2044 72014 2096 72020
rect 2056 71602 2084 72014
rect 2044 71596 2096 71602
rect 2044 71538 2096 71544
rect 1952 70916 2004 70922
rect 1952 70858 2004 70864
rect 1952 70440 2004 70446
rect 1952 70382 2004 70388
rect 1860 68468 1912 68474
rect 1860 68410 1912 68416
rect 1688 68190 1900 68218
rect 1768 68128 1820 68134
rect 1768 68070 1820 68076
rect 1676 67652 1728 67658
rect 1676 67594 1728 67600
rect 1688 67153 1716 67594
rect 1674 67144 1730 67153
rect 1674 67079 1730 67088
rect 1676 67040 1728 67046
rect 1676 66982 1728 66988
rect 1688 60858 1716 66982
rect 1676 60852 1728 60858
rect 1676 60794 1728 60800
rect 1780 58682 1808 68070
rect 1768 58676 1820 58682
rect 1768 58618 1820 58624
rect 1596 58534 1808 58562
rect 1584 58336 1636 58342
rect 1584 58278 1636 58284
rect 1674 58304 1730 58313
rect 1490 58168 1546 58177
rect 1490 58103 1546 58112
rect 1412 58002 1532 58018
rect 1412 57996 1544 58002
rect 1412 57990 1492 57996
rect 1492 57938 1544 57944
rect 1400 57928 1452 57934
rect 1400 57870 1452 57876
rect 1412 57594 1440 57870
rect 1400 57588 1452 57594
rect 1400 57530 1452 57536
rect 1504 57390 1532 57938
rect 1492 57384 1544 57390
rect 1492 57326 1544 57332
rect 1400 57316 1452 57322
rect 1400 57258 1452 57264
rect 1308 56704 1360 56710
rect 1308 56646 1360 56652
rect 1216 53780 1268 53786
rect 1216 53722 1268 53728
rect 1228 52630 1256 53722
rect 1216 52624 1268 52630
rect 1216 52566 1268 52572
rect 1320 51241 1348 56646
rect 1412 56506 1440 57258
rect 1504 56846 1532 57326
rect 1492 56840 1544 56846
rect 1492 56782 1544 56788
rect 1400 56500 1452 56506
rect 1400 56442 1452 56448
rect 1400 56364 1452 56370
rect 1400 56306 1452 56312
rect 1412 55321 1440 56306
rect 1492 56160 1544 56166
rect 1492 56102 1544 56108
rect 1504 55865 1532 56102
rect 1490 55856 1546 55865
rect 1490 55791 1546 55800
rect 1492 55616 1544 55622
rect 1492 55558 1544 55564
rect 1504 55457 1532 55558
rect 1490 55448 1546 55457
rect 1490 55383 1546 55392
rect 1398 55312 1454 55321
rect 1398 55247 1454 55256
rect 1492 55072 1544 55078
rect 1492 55014 1544 55020
rect 1400 54528 1452 54534
rect 1504 54505 1532 55014
rect 1400 54470 1452 54476
rect 1490 54496 1546 54505
rect 1412 53689 1440 54470
rect 1490 54431 1546 54440
rect 1492 53984 1544 53990
rect 1492 53926 1544 53932
rect 1398 53680 1454 53689
rect 1398 53615 1454 53624
rect 1400 53440 1452 53446
rect 1400 53382 1452 53388
rect 1412 51785 1440 53382
rect 1504 52737 1532 53926
rect 1490 52728 1546 52737
rect 1490 52663 1546 52672
rect 1492 52488 1544 52494
rect 1492 52430 1544 52436
rect 1504 51950 1532 52430
rect 1492 51944 1544 51950
rect 1492 51886 1544 51892
rect 1596 51814 1624 58278
rect 1674 58239 1730 58248
rect 1688 57934 1716 58239
rect 1676 57928 1728 57934
rect 1676 57870 1728 57876
rect 1676 57452 1728 57458
rect 1676 57394 1728 57400
rect 1688 57050 1716 57394
rect 1676 57044 1728 57050
rect 1676 56986 1728 56992
rect 1676 56908 1728 56914
rect 1676 56850 1728 56856
rect 1584 51808 1636 51814
rect 1398 51776 1454 51785
rect 1584 51750 1636 51756
rect 1398 51711 1454 51720
rect 1688 51626 1716 56850
rect 1412 51598 1716 51626
rect 1306 51232 1362 51241
rect 1306 51167 1362 51176
rect 1308 51060 1360 51066
rect 1308 51002 1360 51008
rect 1216 50176 1268 50182
rect 1216 50118 1268 50124
rect 1124 49292 1176 49298
rect 1124 49234 1176 49240
rect 1124 49156 1176 49162
rect 1124 49098 1176 49104
rect 1032 47116 1084 47122
rect 1032 47058 1084 47064
rect 1136 47002 1164 49098
rect 1044 46974 1164 47002
rect 940 42764 992 42770
rect 940 42706 992 42712
rect 756 42696 808 42702
rect 1044 42650 1072 46974
rect 1124 46708 1176 46714
rect 1124 46650 1176 46656
rect 756 42638 808 42644
rect 860 42622 1072 42650
rect 860 42514 888 42622
rect 768 42486 888 42514
rect 940 42492 992 42498
rect 664 26444 716 26450
rect 664 26386 716 26392
rect 768 19922 796 42486
rect 940 42434 992 42440
rect 848 42424 900 42430
rect 848 42366 900 42372
rect 756 19916 808 19922
rect 756 19858 808 19864
rect 860 18154 888 42366
rect 952 39030 980 42434
rect 1136 41414 1164 46650
rect 1228 41546 1256 50118
rect 1320 47546 1348 51002
rect 1412 49434 1440 51598
rect 1780 51524 1808 58534
rect 1872 56846 1900 68190
rect 1964 66298 1992 70382
rect 2056 69494 2084 71538
rect 2044 69488 2096 69494
rect 2044 69430 2096 69436
rect 2044 69352 2096 69358
rect 2044 69294 2096 69300
rect 1952 66292 2004 66298
rect 1952 66234 2004 66240
rect 1952 66156 2004 66162
rect 1952 66098 2004 66104
rect 1964 65793 1992 66098
rect 1950 65784 2006 65793
rect 1950 65719 2006 65728
rect 1952 65476 2004 65482
rect 1952 65418 2004 65424
rect 1964 65249 1992 65418
rect 1950 65240 2006 65249
rect 1950 65175 2006 65184
rect 1952 65068 2004 65074
rect 1952 65010 2004 65016
rect 1964 62218 1992 65010
rect 1952 62212 2004 62218
rect 1952 62154 2004 62160
rect 1950 62112 2006 62121
rect 1950 62047 2006 62056
rect 1964 57050 1992 62047
rect 2056 58002 2084 69294
rect 2148 68134 2176 72762
rect 2240 72010 2268 75398
rect 2320 75336 2372 75342
rect 2320 75278 2372 75284
rect 2332 74866 2360 75278
rect 2320 74860 2372 74866
rect 2320 74802 2372 74808
rect 2320 74248 2372 74254
rect 2320 74190 2372 74196
rect 2332 73778 2360 74190
rect 2424 73914 2452 77318
rect 2884 76922 2912 77318
rect 2976 77042 3004 78231
rect 2964 77036 3016 77042
rect 2964 76978 3016 76984
rect 2884 76894 3004 76922
rect 2504 76832 2556 76838
rect 2504 76774 2556 76780
rect 2516 74254 2544 76774
rect 2582 76732 2890 76752
rect 2582 76730 2588 76732
rect 2644 76730 2668 76732
rect 2724 76730 2748 76732
rect 2804 76730 2828 76732
rect 2884 76730 2890 76732
rect 2644 76678 2646 76730
rect 2826 76678 2828 76730
rect 2582 76676 2588 76678
rect 2644 76676 2668 76678
rect 2724 76676 2748 76678
rect 2804 76676 2828 76678
rect 2884 76676 2890 76678
rect 2582 76656 2890 76676
rect 2582 75644 2890 75664
rect 2582 75642 2588 75644
rect 2644 75642 2668 75644
rect 2724 75642 2748 75644
rect 2804 75642 2828 75644
rect 2884 75642 2890 75644
rect 2644 75590 2646 75642
rect 2826 75590 2828 75642
rect 2582 75588 2588 75590
rect 2644 75588 2668 75590
rect 2724 75588 2748 75590
rect 2804 75588 2828 75590
rect 2884 75588 2890 75590
rect 2582 75568 2890 75588
rect 2780 75336 2832 75342
rect 2780 75278 2832 75284
rect 2596 75200 2648 75206
rect 2596 75142 2648 75148
rect 2608 74866 2636 75142
rect 2596 74860 2648 74866
rect 2596 74802 2648 74808
rect 2792 74769 2820 75278
rect 2976 75018 3004 76894
rect 3068 76498 3096 79183
rect 3056 76492 3108 76498
rect 3056 76434 3108 76440
rect 3160 76430 3188 79591
rect 9494 79384 9550 79393
rect 9494 79319 9550 79328
rect 3974 78840 4030 78849
rect 3974 78775 4030 78784
rect 3988 77518 4016 78775
rect 5845 77820 6153 77840
rect 5845 77818 5851 77820
rect 5907 77818 5931 77820
rect 5987 77818 6011 77820
rect 6067 77818 6091 77820
rect 6147 77818 6153 77820
rect 5907 77766 5909 77818
rect 6089 77766 6091 77818
rect 5845 77764 5851 77766
rect 5907 77764 5931 77766
rect 5987 77764 6011 77766
rect 6067 77764 6091 77766
rect 6147 77764 6153 77766
rect 5845 77744 6153 77764
rect 9109 77820 9417 77840
rect 9109 77818 9115 77820
rect 9171 77818 9195 77820
rect 9251 77818 9275 77820
rect 9331 77818 9355 77820
rect 9411 77818 9417 77820
rect 9171 77766 9173 77818
rect 9353 77766 9355 77818
rect 9109 77764 9115 77766
rect 9171 77764 9195 77766
rect 9251 77764 9275 77766
rect 9331 77764 9355 77766
rect 9411 77764 9417 77766
rect 9109 77744 9417 77764
rect 9508 77518 9536 79319
rect 10966 78296 11022 78305
rect 10966 78231 10968 78240
rect 11020 78231 11022 78240
rect 10968 78202 11020 78208
rect 3976 77512 4028 77518
rect 3976 77454 4028 77460
rect 9496 77512 9548 77518
rect 9496 77454 9548 77460
rect 10140 77512 10192 77518
rect 10140 77454 10192 77460
rect 5540 77376 5592 77382
rect 5540 77318 5592 77324
rect 9680 77376 9732 77382
rect 9680 77318 9732 77324
rect 4213 77276 4521 77296
rect 4213 77274 4219 77276
rect 4275 77274 4299 77276
rect 4355 77274 4379 77276
rect 4435 77274 4459 77276
rect 4515 77274 4521 77276
rect 4275 77222 4277 77274
rect 4457 77222 4459 77274
rect 4213 77220 4219 77222
rect 4275 77220 4299 77222
rect 4355 77220 4379 77222
rect 4435 77220 4459 77222
rect 4515 77220 4521 77222
rect 4213 77200 4521 77220
rect 3148 76424 3200 76430
rect 3148 76366 3200 76372
rect 3516 76356 3568 76362
rect 3516 76298 3568 76304
rect 3148 76288 3200 76294
rect 3148 76230 3200 76236
rect 2884 74990 3004 75018
rect 2884 74934 2912 74990
rect 3160 74934 3188 76230
rect 2872 74928 2924 74934
rect 2872 74870 2924 74876
rect 3148 74928 3200 74934
rect 3148 74870 3200 74876
rect 2778 74760 2834 74769
rect 2778 74695 2834 74704
rect 2964 74656 3016 74662
rect 2964 74598 3016 74604
rect 2582 74556 2890 74576
rect 2582 74554 2588 74556
rect 2644 74554 2668 74556
rect 2724 74554 2748 74556
rect 2804 74554 2828 74556
rect 2884 74554 2890 74556
rect 2644 74502 2646 74554
rect 2826 74502 2828 74554
rect 2582 74500 2588 74502
rect 2644 74500 2668 74502
rect 2724 74500 2748 74502
rect 2804 74500 2828 74502
rect 2884 74500 2890 74502
rect 2582 74480 2890 74500
rect 2596 74316 2648 74322
rect 2596 74258 2648 74264
rect 2504 74248 2556 74254
rect 2504 74190 2556 74196
rect 2412 73908 2464 73914
rect 2412 73850 2464 73856
rect 2320 73772 2372 73778
rect 2320 73714 2372 73720
rect 2332 73166 2360 73714
rect 2608 73658 2636 74258
rect 2780 74248 2832 74254
rect 2780 74190 2832 74196
rect 2872 74248 2924 74254
rect 2872 74190 2924 74196
rect 2792 73778 2820 74190
rect 2884 73817 2912 74190
rect 2870 73808 2926 73817
rect 2780 73772 2832 73778
rect 2870 73743 2926 73752
rect 2780 73714 2832 73720
rect 2412 73636 2464 73642
rect 2412 73578 2464 73584
rect 2516 73630 2636 73658
rect 2320 73160 2372 73166
rect 2320 73102 2372 73108
rect 2332 72078 2360 73102
rect 2320 72072 2372 72078
rect 2320 72014 2372 72020
rect 2228 72004 2280 72010
rect 2228 71946 2280 71952
rect 2320 71936 2372 71942
rect 2320 71878 2372 71884
rect 2332 71126 2360 71878
rect 2320 71120 2372 71126
rect 2320 71062 2372 71068
rect 2320 70984 2372 70990
rect 2320 70926 2372 70932
rect 2228 70848 2280 70854
rect 2228 70790 2280 70796
rect 2240 69850 2268 70790
rect 2332 70446 2360 70926
rect 2320 70440 2372 70446
rect 2320 70382 2372 70388
rect 2240 69822 2360 69850
rect 2228 69760 2280 69766
rect 2228 69702 2280 69708
rect 2240 68649 2268 69702
rect 2332 69057 2360 69822
rect 2318 69048 2374 69057
rect 2318 68983 2374 68992
rect 2320 68944 2372 68950
rect 2320 68886 2372 68892
rect 2226 68640 2282 68649
rect 2226 68575 2282 68584
rect 2228 68468 2280 68474
rect 2228 68410 2280 68416
rect 2136 68128 2188 68134
rect 2136 68070 2188 68076
rect 2136 66292 2188 66298
rect 2136 66234 2188 66240
rect 2148 58070 2176 66234
rect 2240 61878 2268 68410
rect 2332 68338 2360 68886
rect 2320 68332 2372 68338
rect 2320 68274 2372 68280
rect 2332 67794 2360 68274
rect 2320 67788 2372 67794
rect 2320 67730 2372 67736
rect 2320 65680 2372 65686
rect 2320 65622 2372 65628
rect 2332 65074 2360 65622
rect 2320 65068 2372 65074
rect 2320 65010 2372 65016
rect 2320 64864 2372 64870
rect 2318 64832 2320 64841
rect 2372 64832 2374 64841
rect 2318 64767 2374 64776
rect 2320 64456 2372 64462
rect 2320 64398 2372 64404
rect 2332 63986 2360 64398
rect 2320 63980 2372 63986
rect 2320 63922 2372 63928
rect 2332 63238 2360 63922
rect 2320 63232 2372 63238
rect 2320 63174 2372 63180
rect 2332 62830 2360 63174
rect 2424 63034 2452 73578
rect 2516 68746 2544 73630
rect 2582 73468 2890 73488
rect 2582 73466 2588 73468
rect 2644 73466 2668 73468
rect 2724 73466 2748 73468
rect 2804 73466 2828 73468
rect 2884 73466 2890 73468
rect 2644 73414 2646 73466
rect 2826 73414 2828 73466
rect 2582 73412 2588 73414
rect 2644 73412 2668 73414
rect 2724 73412 2748 73414
rect 2804 73412 2828 73414
rect 2884 73412 2890 73414
rect 2582 73392 2890 73412
rect 2582 72380 2890 72400
rect 2582 72378 2588 72380
rect 2644 72378 2668 72380
rect 2724 72378 2748 72380
rect 2804 72378 2828 72380
rect 2884 72378 2890 72380
rect 2644 72326 2646 72378
rect 2826 72326 2828 72378
rect 2582 72324 2588 72326
rect 2644 72324 2668 72326
rect 2724 72324 2748 72326
rect 2804 72324 2828 72326
rect 2884 72324 2890 72326
rect 2582 72304 2890 72324
rect 2582 71292 2890 71312
rect 2582 71290 2588 71292
rect 2644 71290 2668 71292
rect 2724 71290 2748 71292
rect 2804 71290 2828 71292
rect 2884 71290 2890 71292
rect 2644 71238 2646 71290
rect 2826 71238 2828 71290
rect 2582 71236 2588 71238
rect 2644 71236 2668 71238
rect 2724 71236 2748 71238
rect 2804 71236 2828 71238
rect 2884 71236 2890 71238
rect 2582 71216 2890 71236
rect 2596 71120 2648 71126
rect 2596 71062 2648 71068
rect 2608 70582 2636 71062
rect 2780 70984 2832 70990
rect 2780 70926 2832 70932
rect 2792 70689 2820 70926
rect 2778 70680 2834 70689
rect 2778 70615 2834 70624
rect 2596 70576 2648 70582
rect 2596 70518 2648 70524
rect 2582 70204 2890 70224
rect 2582 70202 2588 70204
rect 2644 70202 2668 70204
rect 2724 70202 2748 70204
rect 2804 70202 2828 70204
rect 2884 70202 2890 70204
rect 2644 70150 2646 70202
rect 2826 70150 2828 70202
rect 2582 70148 2588 70150
rect 2644 70148 2668 70150
rect 2724 70148 2748 70150
rect 2804 70148 2828 70150
rect 2884 70148 2890 70150
rect 2582 70128 2890 70148
rect 2872 69896 2924 69902
rect 2870 69864 2872 69873
rect 2924 69864 2926 69873
rect 2870 69799 2926 69808
rect 2582 69116 2890 69136
rect 2582 69114 2588 69116
rect 2644 69114 2668 69116
rect 2724 69114 2748 69116
rect 2804 69114 2828 69116
rect 2884 69114 2890 69116
rect 2644 69062 2646 69114
rect 2826 69062 2828 69114
rect 2582 69060 2588 69062
rect 2644 69060 2668 69062
rect 2724 69060 2748 69062
rect 2804 69060 2828 69062
rect 2884 69060 2890 69062
rect 2582 69040 2890 69060
rect 2504 68740 2556 68746
rect 2504 68682 2556 68688
rect 2596 68672 2648 68678
rect 2516 68620 2596 68626
rect 2516 68614 2648 68620
rect 2516 68598 2636 68614
rect 2412 63028 2464 63034
rect 2412 62970 2464 62976
rect 2516 62914 2544 68598
rect 2582 68028 2890 68048
rect 2582 68026 2588 68028
rect 2644 68026 2668 68028
rect 2724 68026 2748 68028
rect 2804 68026 2828 68028
rect 2884 68026 2890 68028
rect 2644 67974 2646 68026
rect 2826 67974 2828 68026
rect 2582 67972 2588 67974
rect 2644 67972 2668 67974
rect 2724 67972 2748 67974
rect 2804 67972 2828 67974
rect 2884 67972 2890 67974
rect 2582 67952 2890 67972
rect 2582 66940 2890 66960
rect 2582 66938 2588 66940
rect 2644 66938 2668 66940
rect 2724 66938 2748 66940
rect 2804 66938 2828 66940
rect 2884 66938 2890 66940
rect 2644 66886 2646 66938
rect 2826 66886 2828 66938
rect 2582 66884 2588 66886
rect 2644 66884 2668 66886
rect 2724 66884 2748 66886
rect 2804 66884 2828 66886
rect 2884 66884 2890 66886
rect 2582 66864 2890 66884
rect 2778 66600 2834 66609
rect 2778 66535 2780 66544
rect 2832 66535 2834 66544
rect 2780 66506 2832 66512
rect 2582 65852 2890 65872
rect 2582 65850 2588 65852
rect 2644 65850 2668 65852
rect 2724 65850 2748 65852
rect 2804 65850 2828 65852
rect 2884 65850 2890 65852
rect 2644 65798 2646 65850
rect 2826 65798 2828 65850
rect 2582 65796 2588 65798
rect 2644 65796 2668 65798
rect 2724 65796 2748 65798
rect 2804 65796 2828 65798
rect 2884 65796 2890 65798
rect 2582 65776 2890 65796
rect 2582 64764 2890 64784
rect 2582 64762 2588 64764
rect 2644 64762 2668 64764
rect 2724 64762 2748 64764
rect 2804 64762 2828 64764
rect 2884 64762 2890 64764
rect 2644 64710 2646 64762
rect 2826 64710 2828 64762
rect 2582 64708 2588 64710
rect 2644 64708 2668 64710
rect 2724 64708 2748 64710
rect 2804 64708 2828 64710
rect 2884 64708 2890 64710
rect 2582 64688 2890 64708
rect 2780 64456 2832 64462
rect 2780 64398 2832 64404
rect 2792 63986 2820 64398
rect 2780 63980 2832 63986
rect 2780 63922 2832 63928
rect 2582 63676 2890 63696
rect 2582 63674 2588 63676
rect 2644 63674 2668 63676
rect 2724 63674 2748 63676
rect 2804 63674 2828 63676
rect 2884 63674 2890 63676
rect 2644 63622 2646 63674
rect 2826 63622 2828 63674
rect 2582 63620 2588 63622
rect 2644 63620 2668 63622
rect 2724 63620 2748 63622
rect 2804 63620 2828 63622
rect 2884 63620 2890 63622
rect 2582 63600 2890 63620
rect 2424 62886 2544 62914
rect 2320 62824 2372 62830
rect 2320 62766 2372 62772
rect 2332 62286 2360 62766
rect 2320 62280 2372 62286
rect 2320 62222 2372 62228
rect 2228 61872 2280 61878
rect 2228 61814 2280 61820
rect 2332 61810 2360 62222
rect 2320 61804 2372 61810
rect 2320 61746 2372 61752
rect 2226 61704 2282 61713
rect 2424 61690 2452 62886
rect 2582 62588 2890 62608
rect 2582 62586 2588 62588
rect 2644 62586 2668 62588
rect 2724 62586 2748 62588
rect 2804 62586 2828 62588
rect 2884 62586 2890 62588
rect 2644 62534 2646 62586
rect 2826 62534 2828 62586
rect 2582 62532 2588 62534
rect 2644 62532 2668 62534
rect 2724 62532 2748 62534
rect 2804 62532 2828 62534
rect 2884 62532 2890 62534
rect 2582 62512 2890 62532
rect 2226 61639 2282 61648
rect 2332 61662 2452 61690
rect 2240 61402 2268 61639
rect 2228 61396 2280 61402
rect 2228 61338 2280 61344
rect 2226 59528 2282 59537
rect 2226 59463 2228 59472
rect 2280 59463 2282 59472
rect 2228 59434 2280 59440
rect 2332 59090 2360 61662
rect 2410 61568 2466 61577
rect 2410 61503 2466 61512
rect 2320 59084 2372 59090
rect 2320 59026 2372 59032
rect 2228 59016 2280 59022
rect 2228 58958 2280 58964
rect 2240 58546 2268 58958
rect 2228 58540 2280 58546
rect 2228 58482 2280 58488
rect 2136 58064 2188 58070
rect 2136 58006 2188 58012
rect 2044 57996 2096 58002
rect 2044 57938 2096 57944
rect 2136 57860 2188 57866
rect 2136 57802 2188 57808
rect 2044 57792 2096 57798
rect 2044 57734 2096 57740
rect 1952 57044 2004 57050
rect 1952 56986 2004 56992
rect 1860 56840 1912 56846
rect 1860 56782 1912 56788
rect 1952 56704 2004 56710
rect 1952 56646 2004 56652
rect 1860 56500 1912 56506
rect 1860 56442 1912 56448
rect 1872 53786 1900 56442
rect 1860 53780 1912 53786
rect 1860 53722 1912 53728
rect 1964 53417 1992 56646
rect 2056 53961 2084 57734
rect 2148 57050 2176 57802
rect 2240 57594 2268 58482
rect 2320 57996 2372 58002
rect 2320 57938 2372 57944
rect 2228 57588 2280 57594
rect 2228 57530 2280 57536
rect 2240 57458 2268 57530
rect 2228 57452 2280 57458
rect 2228 57394 2280 57400
rect 2136 57044 2188 57050
rect 2136 56986 2188 56992
rect 2240 56846 2268 57394
rect 2228 56840 2280 56846
rect 2228 56782 2280 56788
rect 2332 56692 2360 57938
rect 2148 56664 2360 56692
rect 2042 53952 2098 53961
rect 2042 53887 2098 53896
rect 2044 53780 2096 53786
rect 2044 53722 2096 53728
rect 1950 53408 2006 53417
rect 1950 53343 2006 53352
rect 1952 53236 2004 53242
rect 1952 53178 2004 53184
rect 1860 53100 1912 53106
rect 1860 53042 1912 53048
rect 1872 51950 1900 53042
rect 1964 52494 1992 53178
rect 2056 53038 2084 53722
rect 2044 53032 2096 53038
rect 2044 52974 2096 52980
rect 2044 52896 2096 52902
rect 2044 52838 2096 52844
rect 1952 52488 2004 52494
rect 1952 52430 2004 52436
rect 1860 51944 1912 51950
rect 1860 51886 1912 51892
rect 1582 51504 1638 51513
rect 1582 51439 1638 51448
rect 1688 51496 1808 51524
rect 1596 51406 1624 51439
rect 1584 51400 1636 51406
rect 1490 51368 1546 51377
rect 1584 51342 1636 51348
rect 1688 51338 1716 51496
rect 1768 51400 1820 51406
rect 1872 51388 1900 51886
rect 1964 51610 1992 52430
rect 1952 51604 2004 51610
rect 1952 51546 2004 51552
rect 1820 51360 1900 51388
rect 1768 51342 1820 51348
rect 1490 51303 1546 51312
rect 1676 51332 1728 51338
rect 1504 49978 1532 51303
rect 1676 51274 1728 51280
rect 1582 51096 1638 51105
rect 1582 51031 1638 51040
rect 1492 49972 1544 49978
rect 1492 49914 1544 49920
rect 1400 49428 1452 49434
rect 1400 49370 1452 49376
rect 1400 49292 1452 49298
rect 1400 49234 1452 49240
rect 1412 47666 1440 49234
rect 1490 49192 1546 49201
rect 1490 49127 1546 49136
rect 1504 49094 1532 49127
rect 1492 49088 1544 49094
rect 1492 49030 1544 49036
rect 1492 48544 1544 48550
rect 1492 48486 1544 48492
rect 1504 48249 1532 48486
rect 1490 48240 1546 48249
rect 1490 48175 1546 48184
rect 1492 48000 1544 48006
rect 1492 47942 1544 47948
rect 1504 47841 1532 47942
rect 1490 47832 1546 47841
rect 1490 47767 1546 47776
rect 1400 47660 1452 47666
rect 1400 47602 1452 47608
rect 1320 47518 1440 47546
rect 1308 46912 1360 46918
rect 1308 46854 1360 46860
rect 1320 45529 1348 46854
rect 1412 46730 1440 47518
rect 1492 47456 1544 47462
rect 1492 47398 1544 47404
rect 1504 46889 1532 47398
rect 1596 47138 1624 51031
rect 1676 50788 1728 50794
rect 1676 50730 1728 50736
rect 1688 48226 1716 50730
rect 1780 50386 1808 51342
rect 1964 51218 1992 51546
rect 1872 51190 1992 51218
rect 1872 50862 1900 51190
rect 1950 51096 2006 51105
rect 1950 51031 2006 51040
rect 1860 50856 1912 50862
rect 1860 50798 1912 50804
rect 1768 50380 1820 50386
rect 1768 50322 1820 50328
rect 1872 50318 1900 50798
rect 1860 50312 1912 50318
rect 1766 50280 1822 50289
rect 1860 50254 1912 50260
rect 1766 50215 1822 50224
rect 1780 48346 1808 50215
rect 1964 50182 1992 51031
rect 1952 50176 2004 50182
rect 1952 50118 2004 50124
rect 1952 49768 2004 49774
rect 1952 49710 2004 49716
rect 1860 49428 1912 49434
rect 1860 49370 1912 49376
rect 1768 48340 1820 48346
rect 1768 48282 1820 48288
rect 1688 48198 1808 48226
rect 1676 48136 1728 48142
rect 1676 48078 1728 48084
rect 1688 47258 1716 48078
rect 1676 47252 1728 47258
rect 1676 47194 1728 47200
rect 1596 47110 1716 47138
rect 1584 47048 1636 47054
rect 1584 46990 1636 46996
rect 1490 46880 1546 46889
rect 1490 46815 1546 46824
rect 1412 46702 1532 46730
rect 1400 46368 1452 46374
rect 1400 46310 1452 46316
rect 1306 45520 1362 45529
rect 1306 45455 1362 45464
rect 1412 45121 1440 46310
rect 1504 46073 1532 46702
rect 1490 46064 1546 46073
rect 1490 45999 1546 46008
rect 1596 45966 1624 46990
rect 1584 45960 1636 45966
rect 1584 45902 1636 45908
rect 1492 45824 1544 45830
rect 1492 45766 1544 45772
rect 1398 45112 1454 45121
rect 1308 45076 1360 45082
rect 1398 45047 1454 45056
rect 1308 45018 1360 45024
rect 1216 41540 1268 41546
rect 1216 41482 1268 41488
rect 1044 41386 1164 41414
rect 1044 41018 1072 41386
rect 1044 40990 1256 41018
rect 1124 40656 1176 40662
rect 1124 40598 1176 40604
rect 1032 40588 1084 40594
rect 1032 40530 1084 40536
rect 940 39024 992 39030
rect 940 38966 992 38972
rect 848 18148 900 18154
rect 848 18090 900 18096
rect 940 17672 992 17678
rect 940 17614 992 17620
rect 952 16833 980 17614
rect 938 16824 994 16833
rect 938 16759 994 16768
rect 112 11076 164 11082
rect 112 11018 164 11024
rect 1044 9994 1072 40530
rect 1032 9988 1084 9994
rect 1032 9930 1084 9936
rect 1136 5574 1164 40598
rect 1228 5914 1256 40990
rect 1320 40882 1348 45018
rect 1400 44736 1452 44742
rect 1504 44713 1532 45766
rect 1584 45620 1636 45626
rect 1584 45562 1636 45568
rect 1596 44849 1624 45562
rect 1582 44840 1638 44849
rect 1582 44775 1638 44784
rect 1584 44736 1636 44742
rect 1400 44678 1452 44684
rect 1490 44704 1546 44713
rect 1412 42158 1440 44678
rect 1584 44678 1636 44684
rect 1490 44639 1546 44648
rect 1492 44396 1544 44402
rect 1492 44338 1544 44344
rect 1504 43790 1532 44338
rect 1596 44169 1624 44678
rect 1688 44470 1716 47110
rect 1676 44464 1728 44470
rect 1676 44406 1728 44412
rect 1674 44296 1730 44305
rect 1674 44231 1730 44240
rect 1582 44160 1638 44169
rect 1582 44095 1638 44104
rect 1688 43790 1716 44231
rect 1492 43784 1544 43790
rect 1492 43726 1544 43732
rect 1676 43784 1728 43790
rect 1676 43726 1728 43732
rect 1504 43314 1532 43726
rect 1584 43648 1636 43654
rect 1584 43590 1636 43596
rect 1492 43308 1544 43314
rect 1492 43250 1544 43256
rect 1492 42560 1544 42566
rect 1492 42502 1544 42508
rect 1400 42152 1452 42158
rect 1400 42094 1452 42100
rect 1400 42016 1452 42022
rect 1504 41993 1532 42502
rect 1596 42242 1624 43590
rect 1676 42696 1728 42702
rect 1676 42638 1728 42644
rect 1688 42362 1716 42638
rect 1676 42356 1728 42362
rect 1676 42298 1728 42304
rect 1596 42214 1716 42242
rect 1584 42152 1636 42158
rect 1584 42094 1636 42100
rect 1400 41958 1452 41964
rect 1490 41984 1546 41993
rect 1412 41449 1440 41958
rect 1490 41919 1546 41928
rect 1492 41472 1544 41478
rect 1398 41440 1454 41449
rect 1492 41414 1544 41420
rect 1398 41375 1454 41384
rect 1504 41041 1532 41414
rect 1490 41032 1546 41041
rect 1490 40967 1546 40976
rect 1492 40928 1544 40934
rect 1320 40854 1440 40882
rect 1492 40870 1544 40876
rect 1308 40724 1360 40730
rect 1308 40666 1360 40672
rect 1216 5908 1268 5914
rect 1216 5850 1268 5856
rect 1124 5568 1176 5574
rect 1124 5510 1176 5516
rect 1320 5370 1348 40666
rect 1412 40594 1440 40854
rect 1504 40633 1532 40870
rect 1490 40624 1546 40633
rect 1400 40588 1452 40594
rect 1490 40559 1546 40568
rect 1400 40530 1452 40536
rect 1400 40452 1452 40458
rect 1400 40394 1452 40400
rect 1412 38434 1440 40394
rect 1492 40384 1544 40390
rect 1492 40326 1544 40332
rect 1504 40225 1532 40326
rect 1490 40216 1546 40225
rect 1490 40151 1546 40160
rect 1492 39840 1544 39846
rect 1492 39782 1544 39788
rect 1504 39681 1532 39782
rect 1490 39672 1546 39681
rect 1490 39607 1546 39616
rect 1492 39296 1544 39302
rect 1490 39264 1492 39273
rect 1544 39264 1546 39273
rect 1490 39199 1546 39208
rect 1596 38962 1624 42094
rect 1688 40361 1716 42214
rect 1674 40352 1730 40361
rect 1674 40287 1730 40296
rect 1676 40180 1728 40186
rect 1676 40122 1728 40128
rect 1584 38956 1636 38962
rect 1584 38898 1636 38904
rect 1490 38856 1546 38865
rect 1490 38791 1492 38800
rect 1544 38791 1546 38800
rect 1492 38762 1544 38768
rect 1412 38406 1624 38434
rect 1398 38312 1454 38321
rect 1398 38247 1454 38256
rect 1412 38010 1440 38247
rect 1492 38208 1544 38214
rect 1492 38150 1544 38156
rect 1400 38004 1452 38010
rect 1400 37946 1452 37952
rect 1504 37913 1532 38150
rect 1490 37904 1546 37913
rect 1490 37839 1546 37848
rect 1492 37800 1544 37806
rect 1492 37742 1544 37748
rect 1504 37330 1532 37742
rect 1492 37324 1544 37330
rect 1492 37266 1544 37272
rect 1596 37210 1624 38406
rect 1412 37182 1624 37210
rect 1412 36378 1440 37182
rect 1584 37120 1636 37126
rect 1584 37062 1636 37068
rect 1492 36576 1544 36582
rect 1596 36553 1624 37062
rect 1688 36582 1716 40122
rect 1780 36786 1808 48198
rect 1872 44305 1900 49370
rect 1858 44296 1914 44305
rect 1858 44231 1914 44240
rect 1860 44192 1912 44198
rect 1860 44134 1912 44140
rect 1872 40186 1900 44134
rect 1964 41750 1992 49710
rect 1952 41744 2004 41750
rect 1952 41686 2004 41692
rect 1952 41540 2004 41546
rect 1952 41482 2004 41488
rect 1860 40180 1912 40186
rect 1860 40122 1912 40128
rect 1858 40080 1914 40089
rect 1858 40015 1914 40024
rect 1872 37942 1900 40015
rect 1860 37936 1912 37942
rect 1860 37878 1912 37884
rect 1860 37800 1912 37806
rect 1860 37742 1912 37748
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1872 36666 1900 37742
rect 1780 36638 1900 36666
rect 1676 36576 1728 36582
rect 1492 36518 1544 36524
rect 1582 36544 1638 36553
rect 1400 36372 1452 36378
rect 1400 36314 1452 36320
rect 1504 36145 1532 36518
rect 1676 36518 1728 36524
rect 1582 36479 1638 36488
rect 1676 36372 1728 36378
rect 1676 36314 1728 36320
rect 1490 36136 1546 36145
rect 1490 36071 1546 36080
rect 1584 36032 1636 36038
rect 1584 35974 1636 35980
rect 1492 35488 1544 35494
rect 1492 35430 1544 35436
rect 1504 34785 1532 35430
rect 1596 35193 1624 35974
rect 1688 35698 1716 36314
rect 1780 36106 1808 36638
rect 1860 36576 1912 36582
rect 1860 36518 1912 36524
rect 1768 36100 1820 36106
rect 1768 36042 1820 36048
rect 1676 35692 1728 35698
rect 1676 35634 1728 35640
rect 1582 35184 1638 35193
rect 1582 35119 1638 35128
rect 1584 34944 1636 34950
rect 1584 34886 1636 34892
rect 1676 34944 1728 34950
rect 1676 34886 1728 34892
rect 1490 34776 1546 34785
rect 1490 34711 1546 34720
rect 1492 34400 1544 34406
rect 1596 34377 1624 34886
rect 1492 34342 1544 34348
rect 1582 34368 1638 34377
rect 1504 33833 1532 34342
rect 1582 34303 1638 34312
rect 1584 33856 1636 33862
rect 1490 33824 1546 33833
rect 1584 33798 1636 33804
rect 1490 33759 1546 33768
rect 1596 33425 1624 33798
rect 1582 33416 1638 33425
rect 1582 33351 1638 33360
rect 1584 33040 1636 33046
rect 1582 33008 1584 33017
rect 1636 33008 1638 33017
rect 1582 32943 1638 32952
rect 1400 32428 1452 32434
rect 1400 32370 1452 32376
rect 1412 31113 1440 32370
rect 1398 31104 1454 31113
rect 1398 31039 1454 31048
rect 1492 28076 1544 28082
rect 1492 28018 1544 28024
rect 1504 26246 1532 28018
rect 1584 27464 1636 27470
rect 1584 27406 1636 27412
rect 1596 27130 1624 27406
rect 1584 27124 1636 27130
rect 1584 27066 1636 27072
rect 1584 26988 1636 26994
rect 1584 26930 1636 26936
rect 1492 26240 1544 26246
rect 1492 26182 1544 26188
rect 1504 26042 1532 26182
rect 1596 26042 1624 26930
rect 1688 26234 1716 34886
rect 1780 32026 1808 36042
rect 1872 34610 1900 36518
rect 1964 36174 1992 41482
rect 2056 37262 2084 52838
rect 2148 52426 2176 56664
rect 2318 56264 2374 56273
rect 2318 56199 2320 56208
rect 2372 56199 2374 56208
rect 2320 56170 2372 56176
rect 2228 55072 2280 55078
rect 2226 55040 2228 55049
rect 2280 55040 2282 55049
rect 2226 54975 2282 54984
rect 2226 54088 2282 54097
rect 2226 54023 2228 54032
rect 2280 54023 2282 54032
rect 2228 53994 2280 54000
rect 2226 53680 2282 53689
rect 2226 53615 2282 53624
rect 2136 52420 2188 52426
rect 2136 52362 2188 52368
rect 2136 52148 2188 52154
rect 2136 52090 2188 52096
rect 2148 51377 2176 52090
rect 2134 51368 2190 51377
rect 2134 51303 2190 51312
rect 2136 51264 2188 51270
rect 2136 51206 2188 51212
rect 2044 37256 2096 37262
rect 2044 37198 2096 37204
rect 2044 36780 2096 36786
rect 2044 36722 2096 36728
rect 1952 36168 2004 36174
rect 1952 36110 2004 36116
rect 1952 36032 2004 36038
rect 1952 35974 2004 35980
rect 1964 35086 1992 35974
rect 2056 35714 2084 36722
rect 2148 35873 2176 51206
rect 2240 49774 2268 53615
rect 2320 53440 2372 53446
rect 2320 53382 2372 53388
rect 2332 53145 2360 53382
rect 2318 53136 2374 53145
rect 2318 53071 2374 53080
rect 2320 52420 2372 52426
rect 2320 52362 2372 52368
rect 2332 51338 2360 52362
rect 2424 52018 2452 61503
rect 2582 61500 2890 61520
rect 2582 61498 2588 61500
rect 2644 61498 2668 61500
rect 2724 61498 2748 61500
rect 2804 61498 2828 61500
rect 2884 61498 2890 61500
rect 2644 61446 2646 61498
rect 2826 61446 2828 61498
rect 2582 61444 2588 61446
rect 2644 61444 2668 61446
rect 2724 61444 2748 61446
rect 2804 61444 2828 61446
rect 2884 61444 2890 61446
rect 2582 61424 2890 61444
rect 2582 60412 2890 60432
rect 2582 60410 2588 60412
rect 2644 60410 2668 60412
rect 2724 60410 2748 60412
rect 2804 60410 2828 60412
rect 2884 60410 2890 60412
rect 2644 60358 2646 60410
rect 2826 60358 2828 60410
rect 2582 60356 2588 60358
rect 2644 60356 2668 60358
rect 2724 60356 2748 60358
rect 2804 60356 2828 60358
rect 2884 60356 2890 60358
rect 2582 60336 2890 60356
rect 2582 59324 2890 59344
rect 2582 59322 2588 59324
rect 2644 59322 2668 59324
rect 2724 59322 2748 59324
rect 2804 59322 2828 59324
rect 2884 59322 2890 59324
rect 2644 59270 2646 59322
rect 2826 59270 2828 59322
rect 2582 59268 2588 59270
rect 2644 59268 2668 59270
rect 2724 59268 2748 59270
rect 2804 59268 2828 59270
rect 2884 59268 2890 59270
rect 2582 59248 2890 59268
rect 2780 58880 2832 58886
rect 2780 58822 2832 58828
rect 2792 58585 2820 58822
rect 2778 58576 2834 58585
rect 2778 58511 2834 58520
rect 2504 58336 2556 58342
rect 2504 58278 2556 58284
rect 2516 57633 2544 58278
rect 2582 58236 2890 58256
rect 2582 58234 2588 58236
rect 2644 58234 2668 58236
rect 2724 58234 2748 58236
rect 2804 58234 2828 58236
rect 2884 58234 2890 58236
rect 2644 58182 2646 58234
rect 2826 58182 2828 58234
rect 2582 58180 2588 58182
rect 2644 58180 2668 58182
rect 2724 58180 2748 58182
rect 2804 58180 2828 58182
rect 2884 58180 2890 58182
rect 2582 58160 2890 58180
rect 2596 58064 2648 58070
rect 2596 58006 2648 58012
rect 2502 57624 2558 57633
rect 2502 57559 2558 57568
rect 2608 57474 2636 58006
rect 2516 57446 2636 57474
rect 2516 56930 2544 57446
rect 2582 57148 2890 57168
rect 2582 57146 2588 57148
rect 2644 57146 2668 57148
rect 2724 57146 2748 57148
rect 2804 57146 2828 57148
rect 2884 57146 2890 57148
rect 2644 57094 2646 57146
rect 2826 57094 2828 57146
rect 2582 57092 2588 57094
rect 2644 57092 2668 57094
rect 2724 57092 2748 57094
rect 2804 57092 2828 57094
rect 2884 57092 2890 57094
rect 2582 57072 2890 57092
rect 2516 56902 2636 56930
rect 2502 56808 2558 56817
rect 2502 56743 2558 56752
rect 2516 56710 2544 56743
rect 2504 56704 2556 56710
rect 2504 56646 2556 56652
rect 2608 56522 2636 56902
rect 2516 56494 2636 56522
rect 2516 53786 2544 56494
rect 2582 56060 2890 56080
rect 2582 56058 2588 56060
rect 2644 56058 2668 56060
rect 2724 56058 2748 56060
rect 2804 56058 2828 56060
rect 2884 56058 2890 56060
rect 2644 56006 2646 56058
rect 2826 56006 2828 56058
rect 2582 56004 2588 56006
rect 2644 56004 2668 56006
rect 2724 56004 2748 56006
rect 2804 56004 2828 56006
rect 2884 56004 2890 56006
rect 2582 55984 2890 56004
rect 2976 55418 3004 74598
rect 3528 74322 3556 76298
rect 4213 76188 4521 76208
rect 4213 76186 4219 76188
rect 4275 76186 4299 76188
rect 4355 76186 4379 76188
rect 4435 76186 4459 76188
rect 4515 76186 4521 76188
rect 4275 76134 4277 76186
rect 4457 76134 4459 76186
rect 4213 76132 4219 76134
rect 4275 76132 4299 76134
rect 4355 76132 4379 76134
rect 4435 76132 4459 76134
rect 4515 76132 4521 76134
rect 4213 76112 4521 76132
rect 4620 75200 4672 75206
rect 4620 75142 4672 75148
rect 4213 75100 4521 75120
rect 4213 75098 4219 75100
rect 4275 75098 4299 75100
rect 4355 75098 4379 75100
rect 4435 75098 4459 75100
rect 4515 75098 4521 75100
rect 4275 75046 4277 75098
rect 4457 75046 4459 75098
rect 4213 75044 4219 75046
rect 4275 75044 4299 75046
rect 4355 75044 4379 75046
rect 4435 75044 4459 75046
rect 4515 75044 4521 75046
rect 4213 75024 4521 75044
rect 3700 74724 3752 74730
rect 3700 74666 3752 74672
rect 3516 74316 3568 74322
rect 3516 74258 3568 74264
rect 3056 73772 3108 73778
rect 3056 73714 3108 73720
rect 3068 73166 3096 73714
rect 3056 73160 3108 73166
rect 3056 73102 3108 73108
rect 3068 72078 3096 73102
rect 3148 73024 3200 73030
rect 3148 72966 3200 72972
rect 3056 72072 3108 72078
rect 3056 72014 3108 72020
rect 3068 71602 3096 72014
rect 3056 71596 3108 71602
rect 3056 71538 3108 71544
rect 3068 69494 3096 71538
rect 3056 69488 3108 69494
rect 3056 69430 3108 69436
rect 3056 69352 3108 69358
rect 3056 69294 3108 69300
rect 3068 68406 3096 69294
rect 3056 68400 3108 68406
rect 3056 68342 3108 68348
rect 3160 66178 3188 72966
rect 3240 71392 3292 71398
rect 3240 71334 3292 71340
rect 3068 66150 3188 66178
rect 3068 65686 3096 66150
rect 3148 65952 3200 65958
rect 3148 65894 3200 65900
rect 3056 65680 3108 65686
rect 3056 65622 3108 65628
rect 3056 65408 3108 65414
rect 3056 65350 3108 65356
rect 3068 64433 3096 65350
rect 3160 64569 3188 65894
rect 3146 64560 3202 64569
rect 3146 64495 3202 64504
rect 3054 64424 3110 64433
rect 3054 64359 3110 64368
rect 3056 63980 3108 63986
rect 3056 63922 3108 63928
rect 3068 62898 3096 63922
rect 3056 62892 3108 62898
rect 3056 62834 3108 62840
rect 3068 62286 3096 62834
rect 3148 62824 3200 62830
rect 3148 62766 3200 62772
rect 3056 62280 3108 62286
rect 3056 62222 3108 62228
rect 3068 61810 3096 62222
rect 3056 61804 3108 61810
rect 3056 61746 3108 61752
rect 3160 60734 3188 62766
rect 3068 60706 3188 60734
rect 3068 57390 3096 60706
rect 3056 57384 3108 57390
rect 3056 57326 3108 57332
rect 3146 57352 3202 57361
rect 3146 57287 3148 57296
rect 3200 57287 3202 57296
rect 3148 57258 3200 57264
rect 3056 56704 3108 56710
rect 3054 56672 3056 56681
rect 3108 56672 3110 56681
rect 3054 56607 3110 56616
rect 3148 56364 3200 56370
rect 3148 56306 3200 56312
rect 3056 55956 3108 55962
rect 3056 55898 3108 55904
rect 2964 55412 3016 55418
rect 2964 55354 3016 55360
rect 3068 55298 3096 55898
rect 3160 55622 3188 56306
rect 3148 55616 3200 55622
rect 3148 55558 3200 55564
rect 2976 55270 3096 55298
rect 3148 55276 3200 55282
rect 2582 54972 2890 54992
rect 2582 54970 2588 54972
rect 2644 54970 2668 54972
rect 2724 54970 2748 54972
rect 2804 54970 2828 54972
rect 2884 54970 2890 54972
rect 2644 54918 2646 54970
rect 2826 54918 2828 54970
rect 2582 54916 2588 54918
rect 2644 54916 2668 54918
rect 2724 54916 2748 54918
rect 2804 54916 2828 54918
rect 2884 54916 2890 54918
rect 2582 54896 2890 54916
rect 2582 53884 2890 53904
rect 2582 53882 2588 53884
rect 2644 53882 2668 53884
rect 2724 53882 2748 53884
rect 2804 53882 2828 53884
rect 2884 53882 2890 53884
rect 2644 53830 2646 53882
rect 2826 53830 2828 53882
rect 2582 53828 2588 53830
rect 2644 53828 2668 53830
rect 2724 53828 2748 53830
rect 2804 53828 2828 53830
rect 2884 53828 2890 53830
rect 2582 53808 2890 53828
rect 2504 53780 2556 53786
rect 2504 53722 2556 53728
rect 2976 53650 3004 55270
rect 3148 55218 3200 55224
rect 2504 53644 2556 53650
rect 2504 53586 2556 53592
rect 2964 53644 3016 53650
rect 2964 53586 3016 53592
rect 2412 52012 2464 52018
rect 2412 51954 2464 51960
rect 2320 51332 2372 51338
rect 2320 51274 2372 51280
rect 2318 51232 2374 51241
rect 2318 51167 2374 51176
rect 2228 49768 2280 49774
rect 2228 49710 2280 49716
rect 2228 49632 2280 49638
rect 2226 49600 2228 49609
rect 2280 49600 2282 49609
rect 2226 49535 2282 49544
rect 2226 48648 2282 48657
rect 2226 48583 2228 48592
rect 2280 48583 2282 48592
rect 2228 48554 2280 48560
rect 2228 47456 2280 47462
rect 2228 47398 2280 47404
rect 2240 47297 2268 47398
rect 2226 47288 2282 47297
rect 2226 47223 2282 47232
rect 2228 46368 2280 46374
rect 2228 46310 2280 46316
rect 2240 45937 2268 46310
rect 2226 45928 2282 45937
rect 2226 45863 2282 45872
rect 2228 45824 2280 45830
rect 2228 45766 2280 45772
rect 2240 44946 2268 45766
rect 2228 44940 2280 44946
rect 2228 44882 2280 44888
rect 2226 44840 2282 44849
rect 2226 44775 2282 44784
rect 2240 43790 2268 44775
rect 2228 43784 2280 43790
rect 2228 43726 2280 43732
rect 2228 42560 2280 42566
rect 2228 42502 2280 42508
rect 2240 42401 2268 42502
rect 2226 42392 2282 42401
rect 2226 42327 2282 42336
rect 2332 41834 2360 51167
rect 2424 46034 2452 51954
rect 2516 50289 2544 53586
rect 2872 53576 2924 53582
rect 2872 53518 2924 53524
rect 2884 52970 2912 53518
rect 3056 53100 3108 53106
rect 3056 53042 3108 53048
rect 2872 52964 2924 52970
rect 2872 52906 2924 52912
rect 2964 52896 3016 52902
rect 2964 52838 3016 52844
rect 2582 52796 2890 52816
rect 2582 52794 2588 52796
rect 2644 52794 2668 52796
rect 2724 52794 2748 52796
rect 2804 52794 2828 52796
rect 2884 52794 2890 52796
rect 2644 52742 2646 52794
rect 2826 52742 2828 52794
rect 2582 52740 2588 52742
rect 2644 52740 2668 52742
rect 2724 52740 2748 52742
rect 2804 52740 2828 52742
rect 2884 52740 2890 52742
rect 2582 52720 2890 52740
rect 2596 52624 2648 52630
rect 2596 52566 2648 52572
rect 2872 52624 2924 52630
rect 2872 52566 2924 52572
rect 2608 52494 2636 52566
rect 2596 52488 2648 52494
rect 2596 52430 2648 52436
rect 2884 51796 2912 52566
rect 2976 52329 3004 52838
rect 2962 52320 3018 52329
rect 2962 52255 3018 52264
rect 2884 51768 3004 51796
rect 2582 51708 2890 51728
rect 2582 51706 2588 51708
rect 2644 51706 2668 51708
rect 2724 51706 2748 51708
rect 2804 51706 2828 51708
rect 2884 51706 2890 51708
rect 2644 51654 2646 51706
rect 2826 51654 2828 51706
rect 2582 51652 2588 51654
rect 2644 51652 2668 51654
rect 2724 51652 2748 51654
rect 2804 51652 2828 51654
rect 2884 51652 2890 51654
rect 2582 51632 2890 51652
rect 2596 51264 2648 51270
rect 2596 51206 2648 51212
rect 2608 50794 2636 51206
rect 2976 50930 3004 51768
rect 2964 50924 3016 50930
rect 2964 50866 3016 50872
rect 2962 50824 3018 50833
rect 2596 50788 2648 50794
rect 3068 50794 3096 53042
rect 2962 50759 3018 50768
rect 3056 50788 3108 50794
rect 2596 50730 2648 50736
rect 2582 50620 2890 50640
rect 2582 50618 2588 50620
rect 2644 50618 2668 50620
rect 2724 50618 2748 50620
rect 2804 50618 2828 50620
rect 2884 50618 2890 50620
rect 2644 50566 2646 50618
rect 2826 50566 2828 50618
rect 2582 50564 2588 50566
rect 2644 50564 2668 50566
rect 2724 50564 2748 50566
rect 2804 50564 2828 50566
rect 2884 50564 2890 50566
rect 2582 50544 2890 50564
rect 2596 50312 2648 50318
rect 2502 50280 2558 50289
rect 2596 50254 2648 50260
rect 2502 50215 2558 50224
rect 2504 50176 2556 50182
rect 2504 50118 2556 50124
rect 2516 50017 2544 50118
rect 2502 50008 2558 50017
rect 2502 49943 2558 49952
rect 2608 49824 2636 50254
rect 2976 49994 3004 50759
rect 3056 50730 3108 50736
rect 3054 50688 3110 50697
rect 3054 50623 3110 50632
rect 2884 49966 3004 49994
rect 2516 49796 2636 49824
rect 2688 49836 2740 49842
rect 2516 48278 2544 49796
rect 2688 49778 2740 49784
rect 2700 49706 2728 49778
rect 2884 49706 2912 49966
rect 2964 49836 3016 49842
rect 2964 49778 3016 49784
rect 2688 49700 2740 49706
rect 2688 49642 2740 49648
rect 2872 49700 2924 49706
rect 2872 49642 2924 49648
rect 2582 49532 2890 49552
rect 2582 49530 2588 49532
rect 2644 49530 2668 49532
rect 2724 49530 2748 49532
rect 2804 49530 2828 49532
rect 2884 49530 2890 49532
rect 2644 49478 2646 49530
rect 2826 49478 2828 49530
rect 2582 49476 2588 49478
rect 2644 49476 2668 49478
rect 2724 49476 2748 49478
rect 2804 49476 2828 49478
rect 2884 49476 2890 49478
rect 2582 49456 2890 49476
rect 2780 49292 2832 49298
rect 2780 49234 2832 49240
rect 2792 48822 2820 49234
rect 2976 49230 3004 49778
rect 2964 49224 3016 49230
rect 2964 49166 3016 49172
rect 2872 49156 2924 49162
rect 2872 49098 2924 49104
rect 2780 48816 2832 48822
rect 2780 48758 2832 48764
rect 2884 48634 2912 49098
rect 2884 48606 3004 48634
rect 2582 48444 2890 48464
rect 2582 48442 2588 48444
rect 2644 48442 2668 48444
rect 2724 48442 2748 48444
rect 2804 48442 2828 48444
rect 2884 48442 2890 48444
rect 2644 48390 2646 48442
rect 2826 48390 2828 48442
rect 2582 48388 2588 48390
rect 2644 48388 2668 48390
rect 2724 48388 2748 48390
rect 2804 48388 2828 48390
rect 2884 48388 2890 48390
rect 2582 48368 2890 48388
rect 2504 48272 2556 48278
rect 2504 48214 2556 48220
rect 2872 48068 2924 48074
rect 2872 48010 2924 48016
rect 2780 48000 2832 48006
rect 2780 47942 2832 47948
rect 2792 47666 2820 47942
rect 2884 47705 2912 48010
rect 2976 47734 3004 48606
rect 2964 47728 3016 47734
rect 2870 47696 2926 47705
rect 2780 47660 2832 47666
rect 2964 47670 3016 47676
rect 2870 47631 2872 47640
rect 2780 47602 2832 47608
rect 2924 47631 2926 47640
rect 2872 47602 2924 47608
rect 2582 47356 2890 47376
rect 2582 47354 2588 47356
rect 2644 47354 2668 47356
rect 2724 47354 2748 47356
rect 2804 47354 2828 47356
rect 2884 47354 2890 47356
rect 2644 47302 2646 47354
rect 2826 47302 2828 47354
rect 2582 47300 2588 47302
rect 2644 47300 2668 47302
rect 2724 47300 2748 47302
rect 2804 47300 2828 47302
rect 2884 47300 2890 47302
rect 2582 47280 2890 47300
rect 2964 46980 3016 46986
rect 2964 46922 3016 46928
rect 2780 46912 2832 46918
rect 2502 46880 2558 46889
rect 2780 46854 2832 46860
rect 2502 46815 2558 46824
rect 2412 46028 2464 46034
rect 2412 45970 2464 45976
rect 2412 45416 2464 45422
rect 2412 45358 2464 45364
rect 2424 44878 2452 45358
rect 2412 44872 2464 44878
rect 2412 44814 2464 44820
rect 2424 44402 2452 44814
rect 2516 44470 2544 46815
rect 2792 46578 2820 46854
rect 2780 46572 2832 46578
rect 2780 46514 2832 46520
rect 2582 46268 2890 46288
rect 2582 46266 2588 46268
rect 2644 46266 2668 46268
rect 2724 46266 2748 46268
rect 2804 46266 2828 46268
rect 2884 46266 2890 46268
rect 2644 46214 2646 46266
rect 2826 46214 2828 46266
rect 2582 46212 2588 46214
rect 2644 46212 2668 46214
rect 2724 46212 2748 46214
rect 2804 46212 2828 46214
rect 2884 46212 2890 46214
rect 2582 46192 2890 46212
rect 2582 45180 2890 45200
rect 2582 45178 2588 45180
rect 2644 45178 2668 45180
rect 2724 45178 2748 45180
rect 2804 45178 2828 45180
rect 2884 45178 2890 45180
rect 2644 45126 2646 45178
rect 2826 45126 2828 45178
rect 2582 45124 2588 45126
rect 2644 45124 2668 45126
rect 2724 45124 2748 45126
rect 2804 45124 2828 45126
rect 2884 45124 2890 45126
rect 2582 45104 2890 45124
rect 2976 45082 3004 46922
rect 3068 46578 3096 50623
rect 3056 46572 3108 46578
rect 3056 46514 3108 46520
rect 3054 46472 3110 46481
rect 3054 46407 3056 46416
rect 3108 46407 3110 46416
rect 3056 46378 3108 46384
rect 3056 46164 3108 46170
rect 3056 46106 3108 46112
rect 2964 45076 3016 45082
rect 2964 45018 3016 45024
rect 2596 44940 2648 44946
rect 2596 44882 2648 44888
rect 2608 44538 2636 44882
rect 2596 44532 2648 44538
rect 2596 44474 2648 44480
rect 2504 44464 2556 44470
rect 2504 44406 2556 44412
rect 2608 44402 2636 44474
rect 2412 44396 2464 44402
rect 2412 44338 2464 44344
rect 2596 44396 2648 44402
rect 2596 44338 2648 44344
rect 2424 44282 2452 44338
rect 2424 44266 2544 44282
rect 2424 44260 2556 44266
rect 2424 44254 2504 44260
rect 2504 44202 2556 44208
rect 2412 44192 2464 44198
rect 2412 44134 2464 44140
rect 2240 41806 2360 41834
rect 2240 38418 2268 41806
rect 2320 41744 2372 41750
rect 2320 41686 2372 41692
rect 2228 38412 2280 38418
rect 2228 38354 2280 38360
rect 2228 38276 2280 38282
rect 2228 38218 2280 38224
rect 2240 36718 2268 38218
rect 2332 37942 2360 41686
rect 2424 41414 2452 44134
rect 2516 43858 2544 44202
rect 2582 44092 2890 44112
rect 2582 44090 2588 44092
rect 2644 44090 2668 44092
rect 2724 44090 2748 44092
rect 2804 44090 2828 44092
rect 2884 44090 2890 44092
rect 2644 44038 2646 44090
rect 2826 44038 2828 44090
rect 2582 44036 2588 44038
rect 2644 44036 2668 44038
rect 2724 44036 2748 44038
rect 2804 44036 2828 44038
rect 2884 44036 2890 44038
rect 2582 44016 2890 44036
rect 2504 43852 2556 43858
rect 2504 43794 2556 43800
rect 2516 43314 2544 43794
rect 2780 43648 2832 43654
rect 2780 43590 2832 43596
rect 2792 43353 2820 43590
rect 2778 43344 2834 43353
rect 2504 43308 2556 43314
rect 2778 43279 2834 43288
rect 2504 43250 2556 43256
rect 2504 43104 2556 43110
rect 2504 43046 2556 43052
rect 2516 42809 2544 43046
rect 2582 43004 2890 43024
rect 2582 43002 2588 43004
rect 2644 43002 2668 43004
rect 2724 43002 2748 43004
rect 2804 43002 2828 43004
rect 2884 43002 2890 43004
rect 2644 42950 2646 43002
rect 2826 42950 2828 43002
rect 2582 42948 2588 42950
rect 2644 42948 2668 42950
rect 2724 42948 2748 42950
rect 2804 42948 2828 42950
rect 2884 42948 2890 42950
rect 2582 42928 2890 42948
rect 2502 42800 2558 42809
rect 2502 42735 2558 42744
rect 2582 41916 2890 41936
rect 2582 41914 2588 41916
rect 2644 41914 2668 41916
rect 2724 41914 2748 41916
rect 2804 41914 2828 41916
rect 2884 41914 2890 41916
rect 2644 41862 2646 41914
rect 2826 41862 2828 41914
rect 2582 41860 2588 41862
rect 2644 41860 2668 41862
rect 2724 41860 2748 41862
rect 2804 41860 2828 41862
rect 2884 41860 2890 41862
rect 2582 41840 2890 41860
rect 2424 41386 2544 41414
rect 2516 40458 2544 41386
rect 2582 40828 2890 40848
rect 2582 40826 2588 40828
rect 2644 40826 2668 40828
rect 2724 40826 2748 40828
rect 2804 40826 2828 40828
rect 2884 40826 2890 40828
rect 2644 40774 2646 40826
rect 2826 40774 2828 40826
rect 2582 40772 2588 40774
rect 2644 40772 2668 40774
rect 2724 40772 2748 40774
rect 2804 40772 2828 40774
rect 2884 40772 2890 40774
rect 2582 40752 2890 40772
rect 2504 40452 2556 40458
rect 2504 40394 2556 40400
rect 2412 40384 2464 40390
rect 2412 40326 2464 40332
rect 2424 40118 2452 40326
rect 2412 40112 2464 40118
rect 2412 40054 2464 40060
rect 2504 40044 2556 40050
rect 2504 39986 2556 39992
rect 2516 39438 2544 39986
rect 2582 39740 2890 39760
rect 2582 39738 2588 39740
rect 2644 39738 2668 39740
rect 2724 39738 2748 39740
rect 2804 39738 2828 39740
rect 2884 39738 2890 39740
rect 2644 39686 2646 39738
rect 2826 39686 2828 39738
rect 2582 39684 2588 39686
rect 2644 39684 2668 39686
rect 2724 39684 2748 39686
rect 2804 39684 2828 39686
rect 2884 39684 2890 39686
rect 2582 39664 2890 39684
rect 2504 39432 2556 39438
rect 2504 39374 2556 39380
rect 2964 39432 3016 39438
rect 2964 39374 3016 39380
rect 2412 39024 2464 39030
rect 2412 38966 2464 38972
rect 2320 37936 2372 37942
rect 2320 37878 2372 37884
rect 2424 37194 2452 38966
rect 2516 38962 2544 39374
rect 2504 38956 2556 38962
rect 2504 38898 2556 38904
rect 2516 38350 2544 38898
rect 2976 38758 3004 39374
rect 2964 38752 3016 38758
rect 2964 38694 3016 38700
rect 2582 38652 2890 38672
rect 2582 38650 2588 38652
rect 2644 38650 2668 38652
rect 2724 38650 2748 38652
rect 2804 38650 2828 38652
rect 2884 38650 2890 38652
rect 2644 38598 2646 38650
rect 2826 38598 2828 38650
rect 2582 38596 2588 38598
rect 2644 38596 2668 38598
rect 2724 38596 2748 38598
rect 2804 38596 2828 38598
rect 2884 38596 2890 38598
rect 2582 38576 2890 38596
rect 2504 38344 2556 38350
rect 2504 38286 2556 38292
rect 2516 37874 2544 38286
rect 2504 37868 2556 37874
rect 2504 37810 2556 37816
rect 2412 37188 2464 37194
rect 2412 37130 2464 37136
rect 2320 37120 2372 37126
rect 2320 37062 2372 37068
rect 2332 36961 2360 37062
rect 2318 36952 2374 36961
rect 2424 36922 2452 37130
rect 2318 36887 2374 36896
rect 2412 36916 2464 36922
rect 2412 36858 2464 36864
rect 2318 36816 2374 36825
rect 2318 36751 2374 36760
rect 2412 36780 2464 36786
rect 2228 36712 2280 36718
rect 2228 36654 2280 36660
rect 2240 36378 2268 36654
rect 2228 36372 2280 36378
rect 2228 36314 2280 36320
rect 2228 36168 2280 36174
rect 2228 36110 2280 36116
rect 2134 35864 2190 35873
rect 2134 35799 2190 35808
rect 2056 35686 2176 35714
rect 2044 35624 2096 35630
rect 2044 35566 2096 35572
rect 1952 35080 2004 35086
rect 1952 35022 2004 35028
rect 1860 34604 1912 34610
rect 1860 34546 1912 34552
rect 2056 33998 2084 35566
rect 2044 33992 2096 33998
rect 2044 33934 2096 33940
rect 2044 33516 2096 33522
rect 2044 33458 2096 33464
rect 1860 33448 1912 33454
rect 1860 33390 1912 33396
rect 1768 32020 1820 32026
rect 1768 31962 1820 31968
rect 1872 31754 1900 33390
rect 2056 32026 2084 33458
rect 2044 32020 2096 32026
rect 2044 31962 2096 31968
rect 1860 31748 1912 31754
rect 1860 31690 1912 31696
rect 1872 30938 1900 31690
rect 1860 30932 1912 30938
rect 1860 30874 1912 30880
rect 2148 30870 2176 35686
rect 2240 30938 2268 36110
rect 2332 35714 2360 36751
rect 2412 36722 2464 36728
rect 2424 35834 2452 36722
rect 2516 35834 2544 37810
rect 2582 37564 2890 37584
rect 2582 37562 2588 37564
rect 2644 37562 2668 37564
rect 2724 37562 2748 37564
rect 2804 37562 2828 37564
rect 2884 37562 2890 37564
rect 2644 37510 2646 37562
rect 2826 37510 2828 37562
rect 2582 37508 2588 37510
rect 2644 37508 2668 37510
rect 2724 37508 2748 37510
rect 2804 37508 2828 37510
rect 2884 37508 2890 37510
rect 2582 37488 2890 37508
rect 2976 37262 3004 38694
rect 2964 37256 3016 37262
rect 2964 37198 3016 37204
rect 2964 37120 3016 37126
rect 2964 37062 3016 37068
rect 2582 36476 2890 36496
rect 2582 36474 2588 36476
rect 2644 36474 2668 36476
rect 2724 36474 2748 36476
rect 2804 36474 2828 36476
rect 2884 36474 2890 36476
rect 2644 36422 2646 36474
rect 2826 36422 2828 36474
rect 2582 36420 2588 36422
rect 2644 36420 2668 36422
rect 2724 36420 2748 36422
rect 2804 36420 2828 36422
rect 2884 36420 2890 36422
rect 2582 36400 2890 36420
rect 2594 35864 2650 35873
rect 2412 35828 2464 35834
rect 2412 35770 2464 35776
rect 2504 35828 2556 35834
rect 2594 35799 2650 35808
rect 2504 35770 2556 35776
rect 2332 35686 2544 35714
rect 2608 35698 2636 35799
rect 2318 35592 2374 35601
rect 2318 35527 2320 35536
rect 2372 35527 2374 35536
rect 2320 35498 2372 35504
rect 2320 33992 2372 33998
rect 2320 33934 2372 33940
rect 2412 33992 2464 33998
rect 2412 33934 2464 33940
rect 2332 33522 2360 33934
rect 2424 33590 2452 33934
rect 2412 33584 2464 33590
rect 2412 33526 2464 33532
rect 2320 33516 2372 33522
rect 2320 33458 2372 33464
rect 2332 32910 2360 33458
rect 2320 32904 2372 32910
rect 2320 32846 2372 32852
rect 2424 31482 2452 33526
rect 2516 32978 2544 35686
rect 2596 35692 2648 35698
rect 2596 35634 2648 35640
rect 2582 35388 2890 35408
rect 2582 35386 2588 35388
rect 2644 35386 2668 35388
rect 2724 35386 2748 35388
rect 2804 35386 2828 35388
rect 2884 35386 2890 35388
rect 2644 35334 2646 35386
rect 2826 35334 2828 35386
rect 2582 35332 2588 35334
rect 2644 35332 2668 35334
rect 2724 35332 2748 35334
rect 2804 35332 2828 35334
rect 2884 35332 2890 35334
rect 2582 35312 2890 35332
rect 2582 34300 2890 34320
rect 2582 34298 2588 34300
rect 2644 34298 2668 34300
rect 2724 34298 2748 34300
rect 2804 34298 2828 34300
rect 2884 34298 2890 34300
rect 2644 34246 2646 34298
rect 2826 34246 2828 34298
rect 2582 34244 2588 34246
rect 2644 34244 2668 34246
rect 2724 34244 2748 34246
rect 2804 34244 2828 34246
rect 2884 34244 2890 34246
rect 2582 34224 2890 34244
rect 2872 33856 2924 33862
rect 2872 33798 2924 33804
rect 2884 33658 2912 33798
rect 2872 33652 2924 33658
rect 2872 33594 2924 33600
rect 2582 33212 2890 33232
rect 2582 33210 2588 33212
rect 2644 33210 2668 33212
rect 2724 33210 2748 33212
rect 2804 33210 2828 33212
rect 2884 33210 2890 33212
rect 2644 33158 2646 33210
rect 2826 33158 2828 33210
rect 2582 33156 2588 33158
rect 2644 33156 2668 33158
rect 2724 33156 2748 33158
rect 2804 33156 2828 33158
rect 2884 33156 2890 33158
rect 2582 33136 2890 33156
rect 2504 32972 2556 32978
rect 2504 32914 2556 32920
rect 2780 32836 2832 32842
rect 2780 32778 2832 32784
rect 2504 32428 2556 32434
rect 2504 32370 2556 32376
rect 2412 31476 2464 31482
rect 2412 31418 2464 31424
rect 2516 31346 2544 32370
rect 2792 32366 2820 32778
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2582 32124 2890 32144
rect 2582 32122 2588 32124
rect 2644 32122 2668 32124
rect 2724 32122 2748 32124
rect 2804 32122 2828 32124
rect 2884 32122 2890 32124
rect 2644 32070 2646 32122
rect 2826 32070 2828 32122
rect 2582 32068 2588 32070
rect 2644 32068 2668 32070
rect 2724 32068 2748 32070
rect 2804 32068 2828 32070
rect 2884 32068 2890 32070
rect 2582 32048 2890 32068
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2792 31657 2820 31758
rect 2778 31648 2834 31657
rect 2778 31583 2834 31592
rect 2320 31340 2372 31346
rect 2320 31282 2372 31288
rect 2504 31340 2556 31346
rect 2504 31282 2556 31288
rect 2228 30932 2280 30938
rect 2228 30874 2280 30880
rect 2136 30864 2188 30870
rect 2136 30806 2188 30812
rect 1860 30728 1912 30734
rect 1860 30670 1912 30676
rect 1872 29850 1900 30670
rect 2332 30394 2360 31282
rect 2320 30388 2372 30394
rect 2320 30330 2372 30336
rect 2228 30252 2280 30258
rect 2228 30194 2280 30200
rect 2320 30252 2372 30258
rect 2320 30194 2372 30200
rect 1860 29844 1912 29850
rect 1860 29786 1912 29792
rect 2044 29640 2096 29646
rect 2044 29582 2096 29588
rect 1952 29164 2004 29170
rect 1952 29106 2004 29112
rect 1860 29096 1912 29102
rect 1860 29038 1912 29044
rect 1872 27606 1900 29038
rect 1964 28558 1992 29106
rect 1952 28552 2004 28558
rect 1952 28494 2004 28500
rect 2056 27606 2084 29582
rect 2240 29306 2268 30194
rect 2228 29300 2280 29306
rect 2228 29242 2280 29248
rect 2332 28937 2360 30194
rect 2516 30190 2544 31282
rect 2582 31036 2890 31056
rect 2582 31034 2588 31036
rect 2644 31034 2668 31036
rect 2724 31034 2748 31036
rect 2804 31034 2828 31036
rect 2884 31034 2890 31036
rect 2644 30982 2646 31034
rect 2826 30982 2828 31034
rect 2582 30980 2588 30982
rect 2644 30980 2668 30982
rect 2724 30980 2748 30982
rect 2804 30980 2828 30982
rect 2884 30980 2890 30982
rect 2582 30960 2890 30980
rect 2780 30728 2832 30734
rect 2780 30670 2832 30676
rect 2504 30184 2556 30190
rect 2792 30161 2820 30670
rect 2504 30126 2556 30132
rect 2778 30152 2834 30161
rect 2778 30087 2834 30096
rect 2582 29948 2890 29968
rect 2582 29946 2588 29948
rect 2644 29946 2668 29948
rect 2724 29946 2748 29948
rect 2804 29946 2828 29948
rect 2884 29946 2890 29948
rect 2644 29894 2646 29946
rect 2826 29894 2828 29946
rect 2582 29892 2588 29894
rect 2644 29892 2668 29894
rect 2724 29892 2748 29894
rect 2804 29892 2828 29894
rect 2884 29892 2890 29894
rect 2582 29872 2890 29892
rect 2318 28928 2374 28937
rect 2318 28863 2374 28872
rect 2582 28860 2890 28880
rect 2582 28858 2588 28860
rect 2644 28858 2668 28860
rect 2724 28858 2748 28860
rect 2804 28858 2828 28860
rect 2884 28858 2890 28860
rect 2644 28806 2646 28858
rect 2826 28806 2828 28858
rect 2582 28804 2588 28806
rect 2644 28804 2668 28806
rect 2724 28804 2748 28806
rect 2804 28804 2828 28806
rect 2884 28804 2890 28806
rect 2582 28784 2890 28804
rect 2136 28552 2188 28558
rect 2136 28494 2188 28500
rect 2872 28552 2924 28558
rect 2872 28494 2924 28500
rect 1860 27600 1912 27606
rect 1860 27542 1912 27548
rect 2044 27600 2096 27606
rect 2044 27542 2096 27548
rect 2148 26926 2176 28494
rect 2884 28082 2912 28494
rect 2976 28218 3004 37062
rect 3068 35894 3096 46106
rect 3160 46050 3188 55218
rect 3252 50833 3280 71334
rect 3332 70508 3384 70514
rect 3332 70450 3384 70456
rect 3344 68814 3372 70450
rect 3424 69352 3476 69358
rect 3424 69294 3476 69300
rect 3332 68808 3384 68814
rect 3332 68750 3384 68756
rect 3344 68338 3372 68750
rect 3332 68332 3384 68338
rect 3332 68274 3384 68280
rect 3436 67794 3464 69294
rect 3516 68400 3568 68406
rect 3516 68342 3568 68348
rect 3424 67788 3476 67794
rect 3424 67730 3476 67736
rect 3424 66496 3476 66502
rect 3424 66438 3476 66444
rect 3332 64456 3384 64462
rect 3332 64398 3384 64404
rect 3344 53242 3372 64398
rect 3436 55962 3464 66438
rect 3528 65074 3556 68342
rect 3608 67788 3660 67794
rect 3608 67730 3660 67736
rect 3516 65068 3568 65074
rect 3516 65010 3568 65016
rect 3528 63442 3556 65010
rect 3516 63436 3568 63442
rect 3516 63378 3568 63384
rect 3528 57934 3556 63378
rect 3620 62830 3648 67730
rect 3608 62824 3660 62830
rect 3608 62766 3660 62772
rect 3712 60734 3740 74666
rect 3976 74112 4028 74118
rect 3976 74054 4028 74060
rect 3884 68944 3936 68950
rect 3884 68886 3936 68892
rect 3792 65544 3844 65550
rect 3792 65486 3844 65492
rect 3620 60706 3740 60734
rect 3516 57928 3568 57934
rect 3516 57870 3568 57876
rect 3528 56506 3556 57870
rect 3516 56500 3568 56506
rect 3516 56442 3568 56448
rect 3424 55956 3476 55962
rect 3424 55898 3476 55904
rect 3620 55865 3648 60706
rect 3700 57248 3752 57254
rect 3700 57190 3752 57196
rect 3606 55856 3662 55865
rect 3606 55791 3662 55800
rect 3712 55706 3740 57190
rect 3528 55678 3740 55706
rect 3332 53236 3384 53242
rect 3332 53178 3384 53184
rect 3332 53100 3384 53106
rect 3332 53042 3384 53048
rect 3344 52902 3372 53042
rect 3332 52896 3384 52902
rect 3332 52838 3384 52844
rect 3344 52494 3372 52838
rect 3332 52488 3384 52494
rect 3332 52430 3384 52436
rect 3344 51950 3372 52430
rect 3332 51944 3384 51950
rect 3332 51886 3384 51892
rect 3238 50824 3294 50833
rect 3238 50759 3294 50768
rect 3344 50386 3372 51886
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50425 3464 51002
rect 3422 50416 3478 50425
rect 3332 50380 3384 50386
rect 3422 50351 3478 50360
rect 3332 50322 3384 50328
rect 3240 50312 3292 50318
rect 3240 50254 3292 50260
rect 3330 50280 3386 50289
rect 3252 49434 3280 50254
rect 3330 50215 3386 50224
rect 3240 49428 3292 49434
rect 3240 49370 3292 49376
rect 3238 49328 3294 49337
rect 3238 49263 3294 49272
rect 3252 46170 3280 49263
rect 3344 48006 3372 50215
rect 3424 49768 3476 49774
rect 3424 49710 3476 49716
rect 3332 48000 3384 48006
rect 3332 47942 3384 47948
rect 3332 47796 3384 47802
rect 3332 47738 3384 47744
rect 3344 47138 3372 47738
rect 3436 47258 3464 49710
rect 3424 47252 3476 47258
rect 3424 47194 3476 47200
rect 3344 47110 3464 47138
rect 3240 46164 3292 46170
rect 3240 46106 3292 46112
rect 3160 46034 3372 46050
rect 3160 46028 3384 46034
rect 3160 46022 3332 46028
rect 3332 45970 3384 45976
rect 3148 45960 3200 45966
rect 3148 45902 3200 45908
rect 3240 45960 3292 45966
rect 3240 45902 3292 45908
rect 3160 43314 3188 45902
rect 3148 43308 3200 43314
rect 3148 43250 3200 43256
rect 3146 43208 3202 43217
rect 3146 43143 3202 43152
rect 3160 37126 3188 43143
rect 3252 39506 3280 45902
rect 3332 45552 3384 45558
rect 3332 45494 3384 45500
rect 3240 39500 3292 39506
rect 3240 39442 3292 39448
rect 3240 37664 3292 37670
rect 3240 37606 3292 37612
rect 3252 37369 3280 37606
rect 3238 37360 3294 37369
rect 3238 37295 3294 37304
rect 3148 37120 3200 37126
rect 3148 37062 3200 37068
rect 3068 35866 3188 35894
rect 3056 34604 3108 34610
rect 3056 34546 3108 34552
rect 3068 34202 3096 34546
rect 3056 34196 3108 34202
rect 3056 34138 3108 34144
rect 3056 33992 3108 33998
rect 3056 33934 3108 33940
rect 3068 32473 3096 33934
rect 3160 33658 3188 35866
rect 3344 35834 3372 45494
rect 3436 40730 3464 47110
rect 3528 46186 3556 55678
rect 3700 55616 3752 55622
rect 3700 55558 3752 55564
rect 3608 55412 3660 55418
rect 3608 55354 3660 55360
rect 3620 50833 3648 55354
rect 3712 51882 3740 55558
rect 3804 52698 3832 65486
rect 3896 60734 3924 68886
rect 3988 64530 4016 74054
rect 4213 74012 4521 74032
rect 4213 74010 4219 74012
rect 4275 74010 4299 74012
rect 4355 74010 4379 74012
rect 4435 74010 4459 74012
rect 4515 74010 4521 74012
rect 4275 73958 4277 74010
rect 4457 73958 4459 74010
rect 4213 73956 4219 73958
rect 4275 73956 4299 73958
rect 4355 73956 4379 73958
rect 4435 73956 4459 73958
rect 4515 73956 4521 73958
rect 4213 73936 4521 73956
rect 4213 72924 4521 72944
rect 4213 72922 4219 72924
rect 4275 72922 4299 72924
rect 4355 72922 4379 72924
rect 4435 72922 4459 72924
rect 4515 72922 4521 72924
rect 4275 72870 4277 72922
rect 4457 72870 4459 72922
rect 4213 72868 4219 72870
rect 4275 72868 4299 72870
rect 4355 72868 4379 72870
rect 4435 72868 4459 72870
rect 4515 72868 4521 72870
rect 4213 72848 4521 72868
rect 4213 71836 4521 71856
rect 4213 71834 4219 71836
rect 4275 71834 4299 71836
rect 4355 71834 4379 71836
rect 4435 71834 4459 71836
rect 4515 71834 4521 71836
rect 4275 71782 4277 71834
rect 4457 71782 4459 71834
rect 4213 71780 4219 71782
rect 4275 71780 4299 71782
rect 4355 71780 4379 71782
rect 4435 71780 4459 71782
rect 4515 71780 4521 71782
rect 4213 71760 4521 71780
rect 4213 70748 4521 70768
rect 4213 70746 4219 70748
rect 4275 70746 4299 70748
rect 4355 70746 4379 70748
rect 4435 70746 4459 70748
rect 4515 70746 4521 70748
rect 4275 70694 4277 70746
rect 4457 70694 4459 70746
rect 4213 70692 4219 70694
rect 4275 70692 4299 70694
rect 4355 70692 4379 70694
rect 4435 70692 4459 70694
rect 4515 70692 4521 70694
rect 4213 70672 4521 70692
rect 4213 69660 4521 69680
rect 4213 69658 4219 69660
rect 4275 69658 4299 69660
rect 4355 69658 4379 69660
rect 4435 69658 4459 69660
rect 4515 69658 4521 69660
rect 4275 69606 4277 69658
rect 4457 69606 4459 69658
rect 4213 69604 4219 69606
rect 4275 69604 4299 69606
rect 4355 69604 4379 69606
rect 4435 69604 4459 69606
rect 4515 69604 4521 69606
rect 4213 69584 4521 69604
rect 4213 68572 4521 68592
rect 4213 68570 4219 68572
rect 4275 68570 4299 68572
rect 4355 68570 4379 68572
rect 4435 68570 4459 68572
rect 4515 68570 4521 68572
rect 4275 68518 4277 68570
rect 4457 68518 4459 68570
rect 4213 68516 4219 68518
rect 4275 68516 4299 68518
rect 4355 68516 4379 68518
rect 4435 68516 4459 68518
rect 4515 68516 4521 68518
rect 4213 68496 4521 68516
rect 4632 68406 4660 75142
rect 5552 74934 5580 77318
rect 7477 77276 7785 77296
rect 7477 77274 7483 77276
rect 7539 77274 7563 77276
rect 7619 77274 7643 77276
rect 7699 77274 7723 77276
rect 7779 77274 7785 77276
rect 7539 77222 7541 77274
rect 7721 77222 7723 77274
rect 7477 77220 7483 77222
rect 7539 77220 7563 77222
rect 7619 77220 7643 77222
rect 7699 77220 7723 77222
rect 7779 77220 7785 77222
rect 7477 77200 7785 77220
rect 5845 76732 6153 76752
rect 5845 76730 5851 76732
rect 5907 76730 5931 76732
rect 5987 76730 6011 76732
rect 6067 76730 6091 76732
rect 6147 76730 6153 76732
rect 5907 76678 5909 76730
rect 6089 76678 6091 76730
rect 5845 76676 5851 76678
rect 5907 76676 5931 76678
rect 5987 76676 6011 76678
rect 6067 76676 6091 76678
rect 6147 76676 6153 76678
rect 5845 76656 6153 76676
rect 9109 76732 9417 76752
rect 9109 76730 9115 76732
rect 9171 76730 9195 76732
rect 9251 76730 9275 76732
rect 9331 76730 9355 76732
rect 9411 76730 9417 76732
rect 9171 76678 9173 76730
rect 9353 76678 9355 76730
rect 9109 76676 9115 76678
rect 9171 76676 9195 76678
rect 9251 76676 9275 76678
rect 9331 76676 9355 76678
rect 9411 76676 9417 76678
rect 9109 76656 9417 76676
rect 7477 76188 7785 76208
rect 7477 76186 7483 76188
rect 7539 76186 7563 76188
rect 7619 76186 7643 76188
rect 7699 76186 7723 76188
rect 7779 76186 7785 76188
rect 7539 76134 7541 76186
rect 7721 76134 7723 76186
rect 7477 76132 7483 76134
rect 7539 76132 7563 76134
rect 7619 76132 7643 76134
rect 7699 76132 7723 76134
rect 7779 76132 7785 76134
rect 7477 76112 7785 76132
rect 5845 75644 6153 75664
rect 5845 75642 5851 75644
rect 5907 75642 5931 75644
rect 5987 75642 6011 75644
rect 6067 75642 6091 75644
rect 6147 75642 6153 75644
rect 5907 75590 5909 75642
rect 6089 75590 6091 75642
rect 5845 75588 5851 75590
rect 5907 75588 5931 75590
rect 5987 75588 6011 75590
rect 6067 75588 6091 75590
rect 6147 75588 6153 75590
rect 5845 75568 6153 75588
rect 9109 75644 9417 75664
rect 9109 75642 9115 75644
rect 9171 75642 9195 75644
rect 9251 75642 9275 75644
rect 9331 75642 9355 75644
rect 9411 75642 9417 75644
rect 9171 75590 9173 75642
rect 9353 75590 9355 75642
rect 9109 75588 9115 75590
rect 9171 75588 9195 75590
rect 9251 75588 9275 75590
rect 9331 75588 9355 75590
rect 9411 75588 9417 75590
rect 9109 75568 9417 75588
rect 7477 75100 7785 75120
rect 7477 75098 7483 75100
rect 7539 75098 7563 75100
rect 7619 75098 7643 75100
rect 7699 75098 7723 75100
rect 7779 75098 7785 75100
rect 7539 75046 7541 75098
rect 7721 75046 7723 75098
rect 7477 75044 7483 75046
rect 7539 75044 7563 75046
rect 7619 75044 7643 75046
rect 7699 75044 7723 75046
rect 7779 75044 7785 75046
rect 7477 75024 7785 75044
rect 9692 75002 9720 77318
rect 10152 77217 10180 77454
rect 10138 77208 10194 77217
rect 10138 77143 10194 77152
rect 9956 76832 10008 76838
rect 9956 76774 10008 76780
rect 9772 76288 9824 76294
rect 9772 76230 9824 76236
rect 9680 74996 9732 75002
rect 9680 74938 9732 74944
rect 5540 74928 5592 74934
rect 5540 74870 5592 74876
rect 5172 74860 5224 74866
rect 5172 74802 5224 74808
rect 4988 73568 5040 73574
rect 4988 73510 5040 73516
rect 4712 68808 4764 68814
rect 4712 68750 4764 68756
rect 4620 68400 4672 68406
rect 4620 68342 4672 68348
rect 4724 68338 4752 68750
rect 4344 68332 4396 68338
rect 4344 68274 4396 68280
rect 4712 68332 4764 68338
rect 4712 68274 4764 68280
rect 4356 67930 4384 68274
rect 4344 67924 4396 67930
rect 4344 67866 4396 67872
rect 4712 67652 4764 67658
rect 4712 67594 4764 67600
rect 4213 67484 4521 67504
rect 4213 67482 4219 67484
rect 4275 67482 4299 67484
rect 4355 67482 4379 67484
rect 4435 67482 4459 67484
rect 4515 67482 4521 67484
rect 4275 67430 4277 67482
rect 4457 67430 4459 67482
rect 4213 67428 4219 67430
rect 4275 67428 4299 67430
rect 4355 67428 4379 67430
rect 4435 67428 4459 67430
rect 4515 67428 4521 67430
rect 4213 67408 4521 67428
rect 4213 66396 4521 66416
rect 4213 66394 4219 66396
rect 4275 66394 4299 66396
rect 4355 66394 4379 66396
rect 4435 66394 4459 66396
rect 4515 66394 4521 66396
rect 4275 66342 4277 66394
rect 4457 66342 4459 66394
rect 4213 66340 4219 66342
rect 4275 66340 4299 66342
rect 4355 66340 4379 66342
rect 4435 66340 4459 66342
rect 4515 66340 4521 66342
rect 4213 66320 4521 66340
rect 4068 66156 4120 66162
rect 4068 66098 4120 66104
rect 3976 64524 4028 64530
rect 3976 64466 4028 64472
rect 3976 64320 4028 64326
rect 3976 64262 4028 64268
rect 3988 64025 4016 64262
rect 3974 64016 4030 64025
rect 3974 63951 4030 63960
rect 3976 63232 4028 63238
rect 3976 63174 4028 63180
rect 3988 63073 4016 63174
rect 3974 63064 4030 63073
rect 3974 62999 4030 63008
rect 3896 60706 4016 60734
rect 3884 59152 3936 59158
rect 3884 59094 3936 59100
rect 3896 54874 3924 59094
rect 3884 54868 3936 54874
rect 3884 54810 3936 54816
rect 3988 54777 4016 60706
rect 3974 54768 4030 54777
rect 3974 54703 4030 54712
rect 3976 54664 4028 54670
rect 3976 54606 4028 54612
rect 3792 52692 3844 52698
rect 3792 52634 3844 52640
rect 3884 52624 3936 52630
rect 3884 52566 3936 52572
rect 3700 51876 3752 51882
rect 3700 51818 3752 51824
rect 3792 51604 3844 51610
rect 3792 51546 3844 51552
rect 3700 51536 3752 51542
rect 3804 51513 3832 51546
rect 3700 51478 3752 51484
rect 3790 51504 3846 51513
rect 3606 50824 3662 50833
rect 3606 50759 3662 50768
rect 3712 50674 3740 51478
rect 3790 51439 3846 51448
rect 3792 51400 3844 51406
rect 3792 51342 3844 51348
rect 3620 50646 3740 50674
rect 3620 46322 3648 50646
rect 3804 50538 3832 51342
rect 3896 50946 3924 52566
rect 3988 51542 4016 54606
rect 4080 53786 4108 66098
rect 4213 65308 4521 65328
rect 4213 65306 4219 65308
rect 4275 65306 4299 65308
rect 4355 65306 4379 65308
rect 4435 65306 4459 65308
rect 4515 65306 4521 65308
rect 4275 65254 4277 65306
rect 4457 65254 4459 65306
rect 4213 65252 4219 65254
rect 4275 65252 4299 65254
rect 4355 65252 4379 65254
rect 4435 65252 4459 65254
rect 4515 65252 4521 65254
rect 4213 65232 4521 65252
rect 4213 64220 4521 64240
rect 4213 64218 4219 64220
rect 4275 64218 4299 64220
rect 4355 64218 4379 64220
rect 4435 64218 4459 64220
rect 4515 64218 4521 64220
rect 4275 64166 4277 64218
rect 4457 64166 4459 64218
rect 4213 64164 4219 64166
rect 4275 64164 4299 64166
rect 4355 64164 4379 64166
rect 4435 64164 4459 64166
rect 4515 64164 4521 64166
rect 4213 64144 4521 64164
rect 4213 63132 4521 63152
rect 4213 63130 4219 63132
rect 4275 63130 4299 63132
rect 4355 63130 4379 63132
rect 4435 63130 4459 63132
rect 4515 63130 4521 63132
rect 4275 63078 4277 63130
rect 4457 63078 4459 63130
rect 4213 63076 4219 63078
rect 4275 63076 4299 63078
rect 4355 63076 4379 63078
rect 4435 63076 4459 63078
rect 4515 63076 4521 63078
rect 4213 63056 4521 63076
rect 4620 62416 4672 62422
rect 4620 62358 4672 62364
rect 4213 62044 4521 62064
rect 4213 62042 4219 62044
rect 4275 62042 4299 62044
rect 4355 62042 4379 62044
rect 4435 62042 4459 62044
rect 4515 62042 4521 62044
rect 4275 61990 4277 62042
rect 4457 61990 4459 62042
rect 4213 61988 4219 61990
rect 4275 61988 4299 61990
rect 4355 61988 4379 61990
rect 4435 61988 4459 61990
rect 4515 61988 4521 61990
rect 4213 61968 4521 61988
rect 4213 60956 4521 60976
rect 4213 60954 4219 60956
rect 4275 60954 4299 60956
rect 4355 60954 4379 60956
rect 4435 60954 4459 60956
rect 4515 60954 4521 60956
rect 4275 60902 4277 60954
rect 4457 60902 4459 60954
rect 4213 60900 4219 60902
rect 4275 60900 4299 60902
rect 4355 60900 4379 60902
rect 4435 60900 4459 60902
rect 4515 60900 4521 60902
rect 4213 60880 4521 60900
rect 4213 59868 4521 59888
rect 4213 59866 4219 59868
rect 4275 59866 4299 59868
rect 4355 59866 4379 59868
rect 4435 59866 4459 59868
rect 4515 59866 4521 59868
rect 4275 59814 4277 59866
rect 4457 59814 4459 59866
rect 4213 59812 4219 59814
rect 4275 59812 4299 59814
rect 4355 59812 4379 59814
rect 4435 59812 4459 59814
rect 4515 59812 4521 59814
rect 4213 59792 4521 59812
rect 4213 58780 4521 58800
rect 4213 58778 4219 58780
rect 4275 58778 4299 58780
rect 4355 58778 4379 58780
rect 4435 58778 4459 58780
rect 4515 58778 4521 58780
rect 4275 58726 4277 58778
rect 4457 58726 4459 58778
rect 4213 58724 4219 58726
rect 4275 58724 4299 58726
rect 4355 58724 4379 58726
rect 4435 58724 4459 58726
rect 4515 58724 4521 58726
rect 4213 58704 4521 58724
rect 4213 57692 4521 57712
rect 4213 57690 4219 57692
rect 4275 57690 4299 57692
rect 4355 57690 4379 57692
rect 4435 57690 4459 57692
rect 4515 57690 4521 57692
rect 4275 57638 4277 57690
rect 4457 57638 4459 57690
rect 4213 57636 4219 57638
rect 4275 57636 4299 57638
rect 4355 57636 4379 57638
rect 4435 57636 4459 57638
rect 4515 57636 4521 57638
rect 4213 57616 4521 57636
rect 4213 56604 4521 56624
rect 4213 56602 4219 56604
rect 4275 56602 4299 56604
rect 4355 56602 4379 56604
rect 4435 56602 4459 56604
rect 4515 56602 4521 56604
rect 4275 56550 4277 56602
rect 4457 56550 4459 56602
rect 4213 56548 4219 56550
rect 4275 56548 4299 56550
rect 4355 56548 4379 56550
rect 4435 56548 4459 56550
rect 4515 56548 4521 56550
rect 4213 56528 4521 56548
rect 4213 55516 4521 55536
rect 4213 55514 4219 55516
rect 4275 55514 4299 55516
rect 4355 55514 4379 55516
rect 4435 55514 4459 55516
rect 4515 55514 4521 55516
rect 4275 55462 4277 55514
rect 4457 55462 4459 55514
rect 4213 55460 4219 55462
rect 4275 55460 4299 55462
rect 4355 55460 4379 55462
rect 4435 55460 4459 55462
rect 4515 55460 4521 55462
rect 4213 55440 4521 55460
rect 4213 54428 4521 54448
rect 4213 54426 4219 54428
rect 4275 54426 4299 54428
rect 4355 54426 4379 54428
rect 4435 54426 4459 54428
rect 4515 54426 4521 54428
rect 4275 54374 4277 54426
rect 4457 54374 4459 54426
rect 4213 54372 4219 54374
rect 4275 54372 4299 54374
rect 4355 54372 4379 54374
rect 4435 54372 4459 54374
rect 4515 54372 4521 54374
rect 4213 54352 4521 54372
rect 4068 53780 4120 53786
rect 4068 53722 4120 53728
rect 4213 53340 4521 53360
rect 4213 53338 4219 53340
rect 4275 53338 4299 53340
rect 4355 53338 4379 53340
rect 4435 53338 4459 53340
rect 4515 53338 4521 53340
rect 4275 53286 4277 53338
rect 4457 53286 4459 53338
rect 4213 53284 4219 53286
rect 4275 53284 4299 53286
rect 4355 53284 4379 53286
rect 4435 53284 4459 53286
rect 4515 53284 4521 53286
rect 4213 53264 4521 53284
rect 4068 53236 4120 53242
rect 4068 53178 4120 53184
rect 3976 51536 4028 51542
rect 3976 51478 4028 51484
rect 3976 51264 4028 51270
rect 3976 51206 4028 51212
rect 3988 51097 4016 51206
rect 3974 51088 4030 51097
rect 3974 51023 4030 51032
rect 4080 50980 4108 53178
rect 4632 53106 4660 62358
rect 4724 56710 4752 67594
rect 4896 61192 4948 61198
rect 4896 61134 4948 61140
rect 4804 58540 4856 58546
rect 4804 58482 4856 58488
rect 4712 56704 4764 56710
rect 4712 56646 4764 56652
rect 4816 56273 4844 58482
rect 4802 56264 4858 56273
rect 4802 56199 4858 56208
rect 4712 55616 4764 55622
rect 4712 55558 4764 55564
rect 4620 53100 4672 53106
rect 4620 53042 4672 53048
rect 4620 52488 4672 52494
rect 4620 52430 4672 52436
rect 4213 52252 4521 52272
rect 4213 52250 4219 52252
rect 4275 52250 4299 52252
rect 4355 52250 4379 52252
rect 4435 52250 4459 52252
rect 4515 52250 4521 52252
rect 4275 52198 4277 52250
rect 4457 52198 4459 52250
rect 4213 52196 4219 52198
rect 4275 52196 4299 52198
rect 4355 52196 4379 52198
rect 4435 52196 4459 52198
rect 4515 52196 4521 52198
rect 4213 52176 4521 52196
rect 4213 51164 4521 51184
rect 4213 51162 4219 51164
rect 4275 51162 4299 51164
rect 4355 51162 4379 51164
rect 4435 51162 4459 51164
rect 4515 51162 4521 51164
rect 4275 51110 4277 51162
rect 4457 51110 4459 51162
rect 4213 51108 4219 51110
rect 4275 51108 4299 51110
rect 4355 51108 4379 51110
rect 4435 51108 4459 51110
rect 4515 51108 4521 51110
rect 4213 51088 4521 51108
rect 4080 50952 4200 50980
rect 3896 50918 4016 50946
rect 3884 50856 3936 50862
rect 3884 50798 3936 50804
rect 3712 50510 3832 50538
rect 3712 49978 3740 50510
rect 3896 50386 3924 50798
rect 3792 50380 3844 50386
rect 3792 50322 3844 50328
rect 3884 50380 3936 50386
rect 3884 50322 3936 50328
rect 3700 49972 3752 49978
rect 3700 49914 3752 49920
rect 3700 49700 3752 49706
rect 3700 49642 3752 49648
rect 3712 48906 3740 49642
rect 3804 49298 3832 50322
rect 3896 49774 3924 50322
rect 3884 49768 3936 49774
rect 3884 49710 3936 49716
rect 3792 49292 3844 49298
rect 3792 49234 3844 49240
rect 3884 49224 3936 49230
rect 3884 49166 3936 49172
rect 3712 48878 3832 48906
rect 3700 48748 3752 48754
rect 3700 48690 3752 48696
rect 3712 46714 3740 48690
rect 3700 46708 3752 46714
rect 3700 46650 3752 46656
rect 3620 46294 3740 46322
rect 3528 46158 3648 46186
rect 3516 46028 3568 46034
rect 3516 45970 3568 45976
rect 3528 40746 3556 45970
rect 3620 41414 3648 46158
rect 3712 45966 3740 46294
rect 3700 45960 3752 45966
rect 3700 45902 3752 45908
rect 3804 44878 3832 48878
rect 3896 47705 3924 49166
rect 3882 47696 3938 47705
rect 3882 47631 3938 47640
rect 3896 47054 3924 47631
rect 3884 47048 3936 47054
rect 3884 46990 3936 46996
rect 3896 46646 3924 46990
rect 3884 46640 3936 46646
rect 3884 46582 3936 46588
rect 3988 45490 4016 50918
rect 4172 50912 4200 50952
rect 4080 50884 4200 50912
rect 3976 45484 4028 45490
rect 3976 45426 4028 45432
rect 3792 44872 3844 44878
rect 3792 44814 3844 44820
rect 4080 43790 4108 50884
rect 4160 50788 4212 50794
rect 4160 50730 4212 50736
rect 4172 50318 4200 50730
rect 4160 50312 4212 50318
rect 4160 50254 4212 50260
rect 4213 50076 4521 50096
rect 4213 50074 4219 50076
rect 4275 50074 4299 50076
rect 4355 50074 4379 50076
rect 4435 50074 4459 50076
rect 4515 50074 4521 50076
rect 4275 50022 4277 50074
rect 4457 50022 4459 50074
rect 4213 50020 4219 50022
rect 4275 50020 4299 50022
rect 4355 50020 4379 50022
rect 4435 50020 4459 50022
rect 4515 50020 4521 50022
rect 4213 50000 4521 50020
rect 4213 48988 4521 49008
rect 4213 48986 4219 48988
rect 4275 48986 4299 48988
rect 4355 48986 4379 48988
rect 4435 48986 4459 48988
rect 4515 48986 4521 48988
rect 4275 48934 4277 48986
rect 4457 48934 4459 48986
rect 4213 48932 4219 48934
rect 4275 48932 4299 48934
rect 4355 48932 4379 48934
rect 4435 48932 4459 48934
rect 4515 48932 4521 48934
rect 4213 48912 4521 48932
rect 4528 48816 4580 48822
rect 4434 48784 4490 48793
rect 4528 48758 4580 48764
rect 4434 48719 4490 48728
rect 4448 48249 4476 48719
rect 4434 48240 4490 48249
rect 4434 48175 4490 48184
rect 4540 48113 4568 48758
rect 4526 48104 4582 48113
rect 4526 48039 4582 48048
rect 4213 47900 4521 47920
rect 4213 47898 4219 47900
rect 4275 47898 4299 47900
rect 4355 47898 4379 47900
rect 4435 47898 4459 47900
rect 4515 47898 4521 47900
rect 4275 47846 4277 47898
rect 4457 47846 4459 47898
rect 4213 47844 4219 47846
rect 4275 47844 4299 47846
rect 4355 47844 4379 47846
rect 4435 47844 4459 47846
rect 4515 47844 4521 47846
rect 4213 47824 4521 47844
rect 4213 46812 4521 46832
rect 4213 46810 4219 46812
rect 4275 46810 4299 46812
rect 4355 46810 4379 46812
rect 4435 46810 4459 46812
rect 4515 46810 4521 46812
rect 4275 46758 4277 46810
rect 4457 46758 4459 46810
rect 4213 46756 4219 46758
rect 4275 46756 4299 46758
rect 4355 46756 4379 46758
rect 4435 46756 4459 46758
rect 4515 46756 4521 46758
rect 4213 46736 4521 46756
rect 4632 46374 4660 52430
rect 4620 46368 4672 46374
rect 4620 46310 4672 46316
rect 4620 46164 4672 46170
rect 4620 46106 4672 46112
rect 4213 45724 4521 45744
rect 4213 45722 4219 45724
rect 4275 45722 4299 45724
rect 4355 45722 4379 45724
rect 4435 45722 4459 45724
rect 4515 45722 4521 45724
rect 4275 45670 4277 45722
rect 4457 45670 4459 45722
rect 4213 45668 4219 45670
rect 4275 45668 4299 45670
rect 4355 45668 4379 45670
rect 4435 45668 4459 45670
rect 4515 45668 4521 45670
rect 4213 45648 4521 45668
rect 4213 44636 4521 44656
rect 4213 44634 4219 44636
rect 4275 44634 4299 44636
rect 4355 44634 4379 44636
rect 4435 44634 4459 44636
rect 4515 44634 4521 44636
rect 4275 44582 4277 44634
rect 4457 44582 4459 44634
rect 4213 44580 4219 44582
rect 4275 44580 4299 44582
rect 4355 44580 4379 44582
rect 4435 44580 4459 44582
rect 4515 44580 4521 44582
rect 4213 44560 4521 44580
rect 4068 43784 4120 43790
rect 3974 43752 4030 43761
rect 4068 43726 4120 43732
rect 3974 43687 4030 43696
rect 3988 43654 4016 43687
rect 3976 43648 4028 43654
rect 3976 43590 4028 43596
rect 4213 43548 4521 43568
rect 4213 43546 4219 43548
rect 4275 43546 4299 43548
rect 4355 43546 4379 43548
rect 4435 43546 4459 43548
rect 4515 43546 4521 43548
rect 4275 43494 4277 43546
rect 4457 43494 4459 43546
rect 4213 43492 4219 43494
rect 4275 43492 4299 43494
rect 4355 43492 4379 43494
rect 4435 43492 4459 43494
rect 4515 43492 4521 43494
rect 4213 43472 4521 43492
rect 4160 43376 4212 43382
rect 4160 43318 4212 43324
rect 4172 42650 4200 43318
rect 4080 42622 4200 42650
rect 4080 42242 4108 42622
rect 4213 42460 4521 42480
rect 4213 42458 4219 42460
rect 4275 42458 4299 42460
rect 4355 42458 4379 42460
rect 4435 42458 4459 42460
rect 4515 42458 4521 42460
rect 4275 42406 4277 42458
rect 4457 42406 4459 42458
rect 4213 42404 4219 42406
rect 4275 42404 4299 42406
rect 4355 42404 4379 42406
rect 4435 42404 4459 42406
rect 4515 42404 4521 42406
rect 4213 42384 4521 42404
rect 4080 42214 4200 42242
rect 4172 41562 4200 42214
rect 3792 41540 3844 41546
rect 3792 41482 3844 41488
rect 4080 41534 4200 41562
rect 3620 41386 3740 41414
rect 3424 40724 3476 40730
rect 3528 40718 3648 40746
rect 3424 40666 3476 40672
rect 3516 36780 3568 36786
rect 3516 36722 3568 36728
rect 3332 35828 3384 35834
rect 3332 35770 3384 35776
rect 3332 35692 3384 35698
rect 3332 35634 3384 35640
rect 3240 34536 3292 34542
rect 3240 34478 3292 34484
rect 3148 33652 3200 33658
rect 3148 33594 3200 33600
rect 3148 33516 3200 33522
rect 3148 33458 3200 33464
rect 3054 32464 3110 32473
rect 3054 32399 3110 32408
rect 3160 32366 3188 33458
rect 3252 33114 3280 34478
rect 3240 33108 3292 33114
rect 3240 33050 3292 33056
rect 3240 32904 3292 32910
rect 3240 32846 3292 32852
rect 3148 32360 3200 32366
rect 3252 32337 3280 32846
rect 3344 32502 3372 35634
rect 3424 33516 3476 33522
rect 3424 33458 3476 33464
rect 3332 32496 3384 32502
rect 3332 32438 3384 32444
rect 3148 32302 3200 32308
rect 3238 32328 3294 32337
rect 3238 32263 3294 32272
rect 3056 31884 3108 31890
rect 3056 31826 3108 31832
rect 3068 29850 3096 31826
rect 3148 30728 3200 30734
rect 3148 30670 3200 30676
rect 3160 30297 3188 30670
rect 3146 30288 3202 30297
rect 3146 30223 3202 30232
rect 3056 29844 3108 29850
rect 3056 29786 3108 29792
rect 3056 29640 3108 29646
rect 3056 29582 3108 29588
rect 3240 29640 3292 29646
rect 3240 29582 3292 29588
rect 2964 28212 3016 28218
rect 2964 28154 3016 28160
rect 2872 28076 2924 28082
rect 2872 28018 2924 28024
rect 2884 27962 2912 28018
rect 3068 27985 3096 29582
rect 3252 29345 3280 29582
rect 3238 29336 3294 29345
rect 3238 29271 3294 29280
rect 3148 29164 3200 29170
rect 3148 29106 3200 29112
rect 3054 27976 3110 27985
rect 2884 27934 3004 27962
rect 2582 27772 2890 27792
rect 2582 27770 2588 27772
rect 2644 27770 2668 27772
rect 2724 27770 2748 27772
rect 2804 27770 2828 27772
rect 2884 27770 2890 27772
rect 2644 27718 2646 27770
rect 2826 27718 2828 27770
rect 2582 27716 2588 27718
rect 2644 27716 2668 27718
rect 2724 27716 2748 27718
rect 2804 27716 2828 27718
rect 2884 27716 2890 27718
rect 2582 27696 2890 27716
rect 2976 27674 3004 27934
rect 3054 27911 3110 27920
rect 2964 27668 3016 27674
rect 2964 27610 3016 27616
rect 3160 27577 3188 29106
rect 3240 28076 3292 28082
rect 3240 28018 3292 28024
rect 3146 27568 3202 27577
rect 3146 27503 3202 27512
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 2240 27169 2268 27406
rect 2226 27160 2282 27169
rect 2226 27095 2282 27104
rect 2228 26988 2280 26994
rect 2228 26930 2280 26936
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2136 26920 2188 26926
rect 2136 26862 2188 26868
rect 2240 26586 2268 26930
rect 2884 26897 2912 26930
rect 2870 26888 2926 26897
rect 2870 26823 2926 26832
rect 2582 26684 2890 26704
rect 2582 26682 2588 26684
rect 2644 26682 2668 26684
rect 2724 26682 2748 26684
rect 2804 26682 2828 26684
rect 2884 26682 2890 26684
rect 2644 26630 2646 26682
rect 2826 26630 2828 26682
rect 2582 26628 2588 26630
rect 2644 26628 2668 26630
rect 2724 26628 2748 26630
rect 2804 26628 2828 26630
rect 2884 26628 2890 26630
rect 2582 26608 2890 26628
rect 2228 26580 2280 26586
rect 2228 26522 2280 26528
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 2044 26376 2096 26382
rect 2044 26318 2096 26324
rect 1688 26206 1808 26234
rect 1492 26036 1544 26042
rect 1492 25978 1544 25984
rect 1584 26036 1636 26042
rect 1584 25978 1636 25984
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1412 24721 1440 25230
rect 1492 24812 1544 24818
rect 1492 24754 1544 24760
rect 1398 24712 1454 24721
rect 1398 24647 1454 24656
rect 1400 24608 1452 24614
rect 1400 24550 1452 24556
rect 1412 23118 1440 24550
rect 1504 23497 1532 24754
rect 1490 23488 1546 23497
rect 1490 23423 1546 23432
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1490 23080 1546 23089
rect 1490 23015 1546 23024
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 21690 1440 22578
rect 1400 21684 1452 21690
rect 1400 21626 1452 21632
rect 1504 21554 1532 23015
rect 1780 22778 1808 26206
rect 1872 25430 1900 26318
rect 2056 26217 2084 26318
rect 2042 26208 2098 26217
rect 2042 26143 2098 26152
rect 2044 25900 2096 25906
rect 2044 25842 2096 25848
rect 2228 25900 2280 25906
rect 2228 25842 2280 25848
rect 2056 25498 2084 25842
rect 2240 25809 2268 25842
rect 2226 25800 2282 25809
rect 2226 25735 2282 25744
rect 2582 25596 2890 25616
rect 2582 25594 2588 25596
rect 2644 25594 2668 25596
rect 2724 25594 2748 25596
rect 2804 25594 2828 25596
rect 2884 25594 2890 25596
rect 2644 25542 2646 25594
rect 2826 25542 2828 25594
rect 2582 25540 2588 25542
rect 2644 25540 2668 25542
rect 2724 25540 2748 25542
rect 2804 25540 2828 25542
rect 2884 25540 2890 25542
rect 2582 25520 2890 25540
rect 2044 25492 2096 25498
rect 2044 25434 2096 25440
rect 1860 25424 1912 25430
rect 1860 25366 1912 25372
rect 2228 25288 2280 25294
rect 2872 25288 2924 25294
rect 2228 25230 2280 25236
rect 2870 25256 2872 25265
rect 2924 25256 2926 25265
rect 2044 25152 2096 25158
rect 2044 25094 2096 25100
rect 2056 24206 2084 25094
rect 2240 24857 2268 25230
rect 2870 25191 2926 25200
rect 2226 24848 2282 24857
rect 2226 24783 2282 24792
rect 2582 24508 2890 24528
rect 2582 24506 2588 24508
rect 2644 24506 2668 24508
rect 2724 24506 2748 24508
rect 2804 24506 2828 24508
rect 2884 24506 2890 24508
rect 2644 24454 2646 24506
rect 2826 24454 2828 24506
rect 2582 24452 2588 24454
rect 2644 24452 2668 24454
rect 2724 24452 2748 24454
rect 2804 24452 2828 24454
rect 2884 24452 2890 24454
rect 2582 24432 2890 24452
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 2872 24200 2924 24206
rect 2872 24142 2924 24148
rect 2044 24064 2096 24070
rect 2044 24006 2096 24012
rect 2136 24064 2188 24070
rect 2884 24041 2912 24142
rect 2136 24006 2188 24012
rect 2870 24032 2926 24041
rect 2056 23730 2084 24006
rect 2148 23798 2176 24006
rect 2870 23967 2926 23976
rect 2136 23792 2188 23798
rect 2136 23734 2188 23740
rect 2044 23724 2096 23730
rect 2044 23666 2096 23672
rect 2964 23724 3016 23730
rect 2964 23666 3016 23672
rect 2042 23624 2098 23633
rect 2042 23559 2098 23568
rect 2056 23186 2084 23559
rect 2582 23420 2890 23440
rect 2582 23418 2588 23420
rect 2644 23418 2668 23420
rect 2724 23418 2748 23420
rect 2804 23418 2828 23420
rect 2884 23418 2890 23420
rect 2644 23366 2646 23418
rect 2826 23366 2828 23418
rect 2582 23364 2588 23366
rect 2644 23364 2668 23366
rect 2724 23364 2748 23366
rect 2804 23364 2828 23366
rect 2884 23364 2890 23366
rect 2582 23344 2890 23364
rect 2976 23186 3004 23666
rect 3068 23322 3096 27406
rect 3252 26518 3280 28018
rect 3344 27470 3372 32438
rect 3436 31414 3464 33458
rect 3528 32570 3556 36722
rect 3620 35894 3648 40718
rect 3712 37874 3740 41386
rect 3804 40390 3832 41482
rect 4080 41154 4108 41534
rect 4213 41372 4521 41392
rect 4213 41370 4219 41372
rect 4275 41370 4299 41372
rect 4355 41370 4379 41372
rect 4435 41370 4459 41372
rect 4515 41370 4521 41372
rect 4275 41318 4277 41370
rect 4457 41318 4459 41370
rect 4213 41316 4219 41318
rect 4275 41316 4299 41318
rect 4355 41316 4379 41318
rect 4435 41316 4459 41318
rect 4515 41316 4521 41318
rect 4213 41296 4521 41316
rect 4080 41126 4200 41154
rect 3976 40724 4028 40730
rect 3976 40666 4028 40672
rect 3792 40384 3844 40390
rect 3792 40326 3844 40332
rect 3700 37868 3752 37874
rect 3700 37810 3752 37816
rect 3792 37256 3844 37262
rect 3792 37198 3844 37204
rect 3620 35866 3740 35894
rect 3608 35828 3660 35834
rect 3608 35770 3660 35776
rect 3516 32564 3568 32570
rect 3516 32506 3568 32512
rect 3424 31408 3476 31414
rect 3424 31350 3476 31356
rect 3424 31272 3476 31278
rect 3424 31214 3476 31220
rect 3436 29306 3464 31214
rect 3424 29300 3476 29306
rect 3424 29242 3476 29248
rect 3516 29164 3568 29170
rect 3516 29106 3568 29112
rect 3528 28529 3556 29106
rect 3620 28694 3648 35770
rect 3712 34950 3740 35866
rect 3700 34944 3752 34950
rect 3700 34886 3752 34892
rect 3804 30938 3832 37198
rect 3988 35894 4016 40666
rect 4172 40474 4200 41126
rect 4080 40446 4200 40474
rect 4080 40066 4108 40446
rect 4213 40284 4521 40304
rect 4213 40282 4219 40284
rect 4275 40282 4299 40284
rect 4355 40282 4379 40284
rect 4435 40282 4459 40284
rect 4515 40282 4521 40284
rect 4275 40230 4277 40282
rect 4457 40230 4459 40282
rect 4213 40228 4219 40230
rect 4275 40228 4299 40230
rect 4355 40228 4379 40230
rect 4435 40228 4459 40230
rect 4515 40228 4521 40230
rect 4213 40208 4521 40228
rect 4632 40186 4660 46106
rect 4620 40180 4672 40186
rect 4620 40122 4672 40128
rect 4080 40038 4200 40066
rect 4172 39386 4200 40038
rect 4080 39358 4200 39386
rect 4080 38978 4108 39358
rect 4213 39196 4521 39216
rect 4213 39194 4219 39196
rect 4275 39194 4299 39196
rect 4355 39194 4379 39196
rect 4435 39194 4459 39196
rect 4515 39194 4521 39196
rect 4275 39142 4277 39194
rect 4457 39142 4459 39194
rect 4213 39140 4219 39142
rect 4275 39140 4299 39142
rect 4355 39140 4379 39142
rect 4435 39140 4459 39142
rect 4515 39140 4521 39142
rect 4213 39120 4521 39140
rect 4080 38950 4200 38978
rect 4172 38298 4200 38950
rect 4620 38956 4672 38962
rect 4620 38898 4672 38904
rect 4252 38752 4304 38758
rect 4252 38694 4304 38700
rect 4264 38350 4292 38694
rect 4632 38350 4660 38898
rect 4080 38270 4200 38298
rect 4252 38344 4304 38350
rect 4252 38286 4304 38292
rect 4620 38344 4672 38350
rect 4620 38286 4672 38292
rect 4080 38010 4108 38270
rect 4213 38108 4521 38128
rect 4213 38106 4219 38108
rect 4275 38106 4299 38108
rect 4355 38106 4379 38108
rect 4435 38106 4459 38108
rect 4515 38106 4521 38108
rect 4275 38054 4277 38106
rect 4457 38054 4459 38106
rect 4213 38052 4219 38054
rect 4275 38052 4299 38054
rect 4355 38052 4379 38054
rect 4435 38052 4459 38054
rect 4515 38052 4521 38054
rect 4213 38032 4521 38052
rect 4068 38004 4120 38010
rect 4068 37946 4120 37952
rect 4632 37874 4660 38286
rect 4160 37868 4212 37874
rect 4160 37810 4212 37816
rect 4620 37868 4672 37874
rect 4620 37810 4672 37816
rect 4172 37194 4200 37810
rect 4160 37188 4212 37194
rect 4160 37130 4212 37136
rect 4213 37020 4521 37040
rect 4213 37018 4219 37020
rect 4275 37018 4299 37020
rect 4355 37018 4379 37020
rect 4435 37018 4459 37020
rect 4515 37018 4521 37020
rect 4275 36966 4277 37018
rect 4457 36966 4459 37018
rect 4213 36964 4219 36966
rect 4275 36964 4299 36966
rect 4355 36964 4379 36966
rect 4435 36964 4459 36966
rect 4515 36964 4521 36966
rect 4213 36944 4521 36964
rect 4632 36786 4660 37810
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 4632 36174 4660 36722
rect 4620 36168 4672 36174
rect 4620 36110 4672 36116
rect 4213 35932 4521 35952
rect 4213 35930 4219 35932
rect 4275 35930 4299 35932
rect 4355 35930 4379 35932
rect 4435 35930 4459 35932
rect 4515 35930 4521 35932
rect 3988 35866 4108 35894
rect 3792 30932 3844 30938
rect 3792 30874 3844 30880
rect 3976 30728 4028 30734
rect 3974 30696 3976 30705
rect 4028 30696 4030 30705
rect 3974 30631 4030 30640
rect 3792 29096 3844 29102
rect 3792 29038 3844 29044
rect 3608 28688 3660 28694
rect 3608 28630 3660 28636
rect 3804 28558 3832 29038
rect 3700 28552 3752 28558
rect 3514 28520 3570 28529
rect 3700 28494 3752 28500
rect 3792 28552 3844 28558
rect 3792 28494 3844 28500
rect 3514 28455 3570 28464
rect 3712 27470 3740 28494
rect 3332 27464 3384 27470
rect 3332 27406 3384 27412
rect 3700 27464 3752 27470
rect 3700 27406 3752 27412
rect 3976 27464 4028 27470
rect 3976 27406 4028 27412
rect 3712 27062 3740 27406
rect 3700 27056 3752 27062
rect 3700 26998 3752 27004
rect 3988 26994 4016 27406
rect 3976 26988 4028 26994
rect 3976 26930 4028 26936
rect 3240 26512 3292 26518
rect 3240 26454 3292 26460
rect 3792 26376 3844 26382
rect 3792 26318 3844 26324
rect 3240 26308 3292 26314
rect 3240 26250 3292 26256
rect 3252 24818 3280 26250
rect 3804 26246 3832 26318
rect 3792 26240 3844 26246
rect 4080 26234 4108 35866
rect 4275 35878 4277 35930
rect 4457 35878 4459 35930
rect 4213 35876 4219 35878
rect 4275 35876 4299 35878
rect 4355 35876 4379 35878
rect 4435 35876 4459 35878
rect 4515 35876 4521 35878
rect 4213 35856 4521 35876
rect 4632 35154 4660 36110
rect 4620 35148 4672 35154
rect 4620 35090 4672 35096
rect 4213 34844 4521 34864
rect 4213 34842 4219 34844
rect 4275 34842 4299 34844
rect 4355 34842 4379 34844
rect 4435 34842 4459 34844
rect 4515 34842 4521 34844
rect 4275 34790 4277 34842
rect 4457 34790 4459 34842
rect 4213 34788 4219 34790
rect 4275 34788 4299 34790
rect 4355 34788 4379 34790
rect 4435 34788 4459 34790
rect 4515 34788 4521 34790
rect 4213 34768 4521 34788
rect 4213 33756 4521 33776
rect 4213 33754 4219 33756
rect 4275 33754 4299 33756
rect 4355 33754 4379 33756
rect 4435 33754 4459 33756
rect 4515 33754 4521 33756
rect 4275 33702 4277 33754
rect 4457 33702 4459 33754
rect 4213 33700 4219 33702
rect 4275 33700 4299 33702
rect 4355 33700 4379 33702
rect 4435 33700 4459 33702
rect 4515 33700 4521 33702
rect 4213 33680 4521 33700
rect 4252 33516 4304 33522
rect 4252 33458 4304 33464
rect 4528 33516 4580 33522
rect 4528 33458 4580 33464
rect 4264 32910 4292 33458
rect 4540 32910 4568 33458
rect 4252 32904 4304 32910
rect 4252 32846 4304 32852
rect 4528 32904 4580 32910
rect 4580 32852 4660 32858
rect 4528 32846 4660 32852
rect 4540 32830 4660 32846
rect 4213 32668 4521 32688
rect 4213 32666 4219 32668
rect 4275 32666 4299 32668
rect 4355 32666 4379 32668
rect 4435 32666 4459 32668
rect 4515 32666 4521 32668
rect 4275 32614 4277 32666
rect 4457 32614 4459 32666
rect 4213 32612 4219 32614
rect 4275 32612 4299 32614
rect 4355 32612 4379 32614
rect 4435 32612 4459 32614
rect 4515 32612 4521 32614
rect 4213 32592 4521 32612
rect 4632 32434 4660 32830
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 4632 31822 4660 32370
rect 4620 31816 4672 31822
rect 4620 31758 4672 31764
rect 4213 31580 4521 31600
rect 4213 31578 4219 31580
rect 4275 31578 4299 31580
rect 4355 31578 4379 31580
rect 4435 31578 4459 31580
rect 4515 31578 4521 31580
rect 4275 31526 4277 31578
rect 4457 31526 4459 31578
rect 4213 31524 4219 31526
rect 4275 31524 4299 31526
rect 4355 31524 4379 31526
rect 4435 31524 4459 31526
rect 4515 31524 4521 31526
rect 4213 31504 4521 31524
rect 4632 31346 4660 31758
rect 4620 31340 4672 31346
rect 4620 31282 4672 31288
rect 4632 30734 4660 31282
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 4213 30492 4521 30512
rect 4213 30490 4219 30492
rect 4275 30490 4299 30492
rect 4355 30490 4379 30492
rect 4435 30490 4459 30492
rect 4515 30490 4521 30492
rect 4275 30438 4277 30490
rect 4457 30438 4459 30490
rect 4213 30436 4219 30438
rect 4275 30436 4299 30438
rect 4355 30436 4379 30438
rect 4435 30436 4459 30438
rect 4515 30436 4521 30438
rect 4213 30416 4521 30436
rect 4213 29404 4521 29424
rect 4213 29402 4219 29404
rect 4275 29402 4299 29404
rect 4355 29402 4379 29404
rect 4435 29402 4459 29404
rect 4515 29402 4521 29404
rect 4275 29350 4277 29402
rect 4457 29350 4459 29402
rect 4213 29348 4219 29350
rect 4275 29348 4299 29350
rect 4355 29348 4379 29350
rect 4435 29348 4459 29350
rect 4515 29348 4521 29350
rect 4213 29328 4521 29348
rect 4620 28552 4672 28558
rect 4620 28494 4672 28500
rect 4213 28316 4521 28336
rect 4213 28314 4219 28316
rect 4275 28314 4299 28316
rect 4355 28314 4379 28316
rect 4435 28314 4459 28316
rect 4515 28314 4521 28316
rect 4275 28262 4277 28314
rect 4457 28262 4459 28314
rect 4213 28260 4219 28262
rect 4275 28260 4299 28262
rect 4355 28260 4379 28262
rect 4435 28260 4459 28262
rect 4515 28260 4521 28262
rect 4213 28240 4521 28260
rect 4528 28076 4580 28082
rect 4528 28018 4580 28024
rect 4252 28008 4304 28014
rect 4252 27950 4304 27956
rect 4264 27470 4292 27950
rect 4540 27826 4568 28018
rect 4632 28014 4660 28494
rect 4620 28008 4672 28014
rect 4620 27950 4672 27956
rect 4540 27798 4660 27826
rect 4252 27464 4304 27470
rect 4252 27406 4304 27412
rect 4213 27228 4521 27248
rect 4213 27226 4219 27228
rect 4275 27226 4299 27228
rect 4355 27226 4379 27228
rect 4435 27226 4459 27228
rect 4515 27226 4521 27228
rect 4275 27174 4277 27226
rect 4457 27174 4459 27226
rect 4213 27172 4219 27174
rect 4275 27172 4299 27174
rect 4355 27172 4379 27174
rect 4435 27172 4459 27174
rect 4515 27172 4521 27174
rect 4213 27152 4521 27172
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4172 26314 4200 26930
rect 4160 26308 4212 26314
rect 4160 26250 4212 26256
rect 3792 26182 3844 26188
rect 3988 26206 4108 26234
rect 3240 24812 3292 24818
rect 3240 24754 3292 24760
rect 3056 23316 3108 23322
rect 3056 23258 3108 23264
rect 2044 23180 2096 23186
rect 2044 23122 2096 23128
rect 2964 23180 3016 23186
rect 2964 23122 3016 23128
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 2976 22642 3004 23122
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 1688 21894 1716 22578
rect 2582 22332 2890 22352
rect 2582 22330 2588 22332
rect 2644 22330 2668 22332
rect 2724 22330 2748 22332
rect 2804 22330 2828 22332
rect 2884 22330 2890 22332
rect 2644 22278 2646 22330
rect 2826 22278 2828 22330
rect 2582 22276 2588 22278
rect 2644 22276 2668 22278
rect 2724 22276 2748 22278
rect 2804 22276 2828 22278
rect 2884 22276 2890 22278
rect 2582 22256 2890 22276
rect 2976 22234 3004 22578
rect 2964 22228 3016 22234
rect 2964 22170 3016 22176
rect 3068 22030 3096 23258
rect 3148 23112 3200 23118
rect 3148 23054 3200 23060
rect 3160 22030 3188 23054
rect 2044 22024 2096 22030
rect 2044 21966 2096 21972
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 3148 22024 3200 22030
rect 3148 21966 3200 21972
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1688 21622 1716 21830
rect 2056 21729 2084 21966
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 2042 21720 2098 21729
rect 2042 21655 2098 21664
rect 1676 21616 1728 21622
rect 1676 21558 1728 21564
rect 1492 21548 1544 21554
rect 1492 21490 1544 21496
rect 1584 21548 1636 21554
rect 1584 21490 1636 21496
rect 1492 20936 1544 20942
rect 1492 20878 1544 20884
rect 1400 20460 1452 20466
rect 1400 20402 1452 20408
rect 1412 19009 1440 20402
rect 1504 19553 1532 20878
rect 1596 20777 1624 21490
rect 1860 21344 1912 21350
rect 1860 21286 1912 21292
rect 2228 21344 2280 21350
rect 2228 21286 2280 21292
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1582 20768 1638 20777
rect 1582 20703 1638 20712
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1490 19544 1546 19553
rect 1490 19479 1546 19488
rect 1398 19000 1454 19009
rect 1398 18935 1454 18944
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17377 1440 18226
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1398 17368 1454 17377
rect 1398 17303 1454 17312
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 1412 16289 1440 17138
rect 1504 16658 1532 18022
rect 1596 17678 1624 20198
rect 1688 19961 1716 20878
rect 1768 20800 1820 20806
rect 1768 20742 1820 20748
rect 1674 19952 1730 19961
rect 1674 19887 1730 19896
rect 1780 18290 1808 20742
rect 1872 19854 1900 21286
rect 2044 20800 2096 20806
rect 2044 20742 2096 20748
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1872 19378 1900 19654
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 2056 18766 2084 20742
rect 2240 20466 2268 21286
rect 2516 20466 2544 21830
rect 2872 21548 2924 21554
rect 2872 21490 2924 21496
rect 2884 21457 2912 21490
rect 2870 21448 2926 21457
rect 2870 21383 2926 21392
rect 2582 21244 2890 21264
rect 2582 21242 2588 21244
rect 2644 21242 2668 21244
rect 2724 21242 2748 21244
rect 2804 21242 2828 21244
rect 2884 21242 2890 21244
rect 2644 21190 2646 21242
rect 2826 21190 2828 21242
rect 2582 21188 2588 21190
rect 2644 21188 2668 21190
rect 2724 21188 2748 21190
rect 2804 21188 2828 21190
rect 2884 21188 2890 21190
rect 2582 21168 2890 21188
rect 3068 20942 3096 21966
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2412 20392 2464 20398
rect 2412 20334 2464 20340
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 2148 18426 2176 19858
rect 2424 19514 2452 20334
rect 2582 20156 2890 20176
rect 2582 20154 2588 20156
rect 2644 20154 2668 20156
rect 2724 20154 2748 20156
rect 2804 20154 2828 20156
rect 2884 20154 2890 20156
rect 2644 20102 2646 20154
rect 2826 20102 2828 20154
rect 2582 20100 2588 20102
rect 2644 20100 2668 20102
rect 2724 20100 2748 20102
rect 2804 20100 2828 20102
rect 2884 20100 2890 20102
rect 2582 20080 2890 20100
rect 2964 19984 3016 19990
rect 2964 19926 3016 19932
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 2516 19378 2544 19790
rect 2976 19514 3004 19926
rect 3068 19922 3096 20742
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 2504 19372 2556 19378
rect 2504 19314 2556 19320
rect 2516 18766 2544 19314
rect 2964 19236 3016 19242
rect 2964 19178 3016 19184
rect 2582 19068 2890 19088
rect 2582 19066 2588 19068
rect 2644 19066 2668 19068
rect 2724 19066 2748 19068
rect 2804 19066 2828 19068
rect 2884 19066 2890 19068
rect 2644 19014 2646 19066
rect 2826 19014 2828 19066
rect 2582 19012 2588 19014
rect 2644 19012 2668 19014
rect 2724 19012 2748 19014
rect 2804 19012 2828 19014
rect 2884 19012 2890 19014
rect 2582 18992 2890 19012
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 2136 18420 2188 18426
rect 2136 18362 2188 18368
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 2044 18148 2096 18154
rect 2044 18090 2096 18096
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1596 16590 1624 17478
rect 2056 17338 2084 18090
rect 2148 18086 2176 18362
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 2582 17980 2890 18000
rect 2582 17978 2588 17980
rect 2644 17978 2668 17980
rect 2724 17978 2748 17980
rect 2804 17978 2828 17980
rect 2884 17978 2890 17980
rect 2644 17926 2646 17978
rect 2826 17926 2828 17978
rect 2582 17924 2588 17926
rect 2644 17924 2668 17926
rect 2724 17924 2748 17926
rect 2804 17924 2828 17926
rect 2884 17924 2890 17926
rect 2582 17904 2890 17924
rect 2872 17672 2924 17678
rect 2870 17640 2872 17649
rect 2924 17640 2926 17649
rect 2870 17575 2926 17584
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1398 16280 1454 16289
rect 1398 16215 1454 16224
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 14521 1440 15438
rect 1504 15065 1532 16050
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1490 15056 1546 15065
rect 1490 14991 1546 15000
rect 1398 14512 1454 14521
rect 1398 14447 1454 14456
rect 1596 14226 1624 15302
rect 1688 15026 1716 16934
rect 2240 16794 2268 17478
rect 2582 16892 2890 16912
rect 2582 16890 2588 16892
rect 2644 16890 2668 16892
rect 2724 16890 2748 16892
rect 2804 16890 2828 16892
rect 2884 16890 2890 16892
rect 2644 16838 2646 16890
rect 2826 16838 2828 16890
rect 2582 16836 2588 16838
rect 2644 16836 2668 16838
rect 2724 16836 2748 16838
rect 2804 16836 2828 16838
rect 2884 16836 2890 16838
rect 2582 16816 2890 16836
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2136 16448 2188 16454
rect 2136 16390 2188 16396
rect 1952 15972 2004 15978
rect 1952 15914 2004 15920
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1780 14482 1808 14758
rect 1872 14618 1900 15846
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1964 14346 1992 15914
rect 2044 15360 2096 15366
rect 2044 15302 2096 15308
rect 2056 15094 2084 15302
rect 2044 15088 2096 15094
rect 2044 15030 2096 15036
rect 2148 14414 2176 16390
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2240 15881 2268 16050
rect 2226 15872 2282 15881
rect 2226 15807 2282 15816
rect 2582 15804 2890 15824
rect 2582 15802 2588 15804
rect 2644 15802 2668 15804
rect 2724 15802 2748 15804
rect 2804 15802 2828 15804
rect 2884 15802 2890 15804
rect 2644 15750 2646 15802
rect 2826 15750 2828 15802
rect 2582 15748 2588 15750
rect 2644 15748 2668 15750
rect 2724 15748 2748 15750
rect 2804 15748 2828 15750
rect 2884 15748 2890 15750
rect 2582 15728 2890 15748
rect 2228 15496 2280 15502
rect 2226 15464 2228 15473
rect 2280 15464 2282 15473
rect 2226 15399 2282 15408
rect 2582 14716 2890 14736
rect 2582 14714 2588 14716
rect 2644 14714 2668 14716
rect 2724 14714 2748 14716
rect 2804 14714 2828 14716
rect 2884 14714 2890 14716
rect 2644 14662 2646 14714
rect 2826 14662 2828 14714
rect 2582 14660 2588 14662
rect 2644 14660 2668 14662
rect 2724 14660 2748 14662
rect 2804 14660 2828 14662
rect 2884 14660 2890 14662
rect 2582 14640 2890 14660
rect 2412 14544 2464 14550
rect 2412 14486 2464 14492
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 2136 14272 2188 14278
rect 1596 14198 1900 14226
rect 2136 14214 2188 14220
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13161 1440 13874
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1398 13152 1454 13161
rect 1398 13087 1454 13096
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 11801 1440 12786
rect 1504 12345 1532 13262
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 1596 12238 1624 12582
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1688 12170 1716 14010
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1584 12096 1636 12102
rect 1636 12044 1716 12050
rect 1584 12038 1716 12044
rect 1596 12022 1716 12038
rect 1398 11792 1454 11801
rect 1398 11727 1454 11736
rect 1398 11384 1454 11393
rect 1688 11354 1716 12022
rect 1780 11558 1808 13126
rect 1872 12238 1900 14198
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1872 11762 1900 12038
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1398 11319 1454 11328
rect 1676 11348 1728 11354
rect 1412 11150 1440 11319
rect 1676 11290 1728 11296
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 10266 1624 10950
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1688 10130 1716 11290
rect 1872 10674 1900 11698
rect 1964 11626 1992 14010
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 2056 11694 2084 12582
rect 2148 11762 2176 14214
rect 2332 14113 2360 14350
rect 2318 14104 2374 14113
rect 2318 14039 2374 14048
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2240 13705 2268 13874
rect 2226 13696 2282 13705
rect 2226 13631 2282 13640
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2240 12753 2268 12786
rect 2226 12744 2282 12753
rect 2226 12679 2282 12688
rect 2424 11914 2452 14486
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2240 11886 2452 11914
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2044 11688 2096 11694
rect 2240 11642 2268 11886
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 2044 11630 2096 11636
rect 1952 11620 2004 11626
rect 1952 11562 2004 11568
rect 2148 11614 2268 11642
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 2056 10062 2084 11494
rect 2148 11150 2176 11614
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2148 10742 2176 11086
rect 2136 10736 2188 10742
rect 2136 10678 2188 10684
rect 2240 10266 2268 11086
rect 2332 10674 2360 11494
rect 2424 11150 2452 11766
rect 2516 11694 2544 14214
rect 2582 13628 2890 13648
rect 2582 13626 2588 13628
rect 2644 13626 2668 13628
rect 2724 13626 2748 13628
rect 2804 13626 2828 13628
rect 2884 13626 2890 13628
rect 2644 13574 2646 13626
rect 2826 13574 2828 13626
rect 2582 13572 2588 13574
rect 2644 13572 2668 13574
rect 2724 13572 2748 13574
rect 2804 13572 2828 13574
rect 2884 13572 2890 13574
rect 2582 13552 2890 13572
rect 2582 12540 2890 12560
rect 2582 12538 2588 12540
rect 2644 12538 2668 12540
rect 2724 12538 2748 12540
rect 2804 12538 2828 12540
rect 2884 12538 2890 12540
rect 2644 12486 2646 12538
rect 2826 12486 2828 12538
rect 2582 12484 2588 12486
rect 2644 12484 2668 12486
rect 2724 12484 2748 12486
rect 2804 12484 2828 12486
rect 2884 12484 2890 12486
rect 2582 12464 2890 12484
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11354 2544 11494
rect 2582 11452 2890 11472
rect 2582 11450 2588 11452
rect 2644 11450 2668 11452
rect 2724 11450 2748 11452
rect 2804 11450 2828 11452
rect 2884 11450 2890 11452
rect 2644 11398 2646 11450
rect 2826 11398 2828 11450
rect 2582 11396 2588 11398
rect 2644 11396 2668 11398
rect 2724 11396 2748 11398
rect 2804 11396 2828 11398
rect 2884 11396 2890 11398
rect 2582 11376 2890 11396
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2976 11218 3004 19178
rect 3068 18766 3096 19654
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 3068 18222 3096 18702
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 3160 18154 3188 19790
rect 3148 18148 3200 18154
rect 3148 18090 3200 18096
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 3068 11150 3096 18022
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2582 10364 2890 10384
rect 2582 10362 2588 10364
rect 2644 10362 2668 10364
rect 2724 10362 2748 10364
rect 2804 10362 2828 10364
rect 2884 10362 2890 10364
rect 2644 10310 2646 10362
rect 2826 10310 2828 10362
rect 2582 10308 2588 10310
rect 2644 10308 2668 10310
rect 2724 10308 2748 10310
rect 2804 10308 2828 10310
rect 2884 10308 2890 10310
rect 2582 10288 2890 10308
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2240 6390 2268 9930
rect 2582 9276 2890 9296
rect 2582 9274 2588 9276
rect 2644 9274 2668 9276
rect 2724 9274 2748 9276
rect 2804 9274 2828 9276
rect 2884 9274 2890 9276
rect 2644 9222 2646 9274
rect 2826 9222 2828 9274
rect 2582 9220 2588 9222
rect 2644 9220 2668 9222
rect 2724 9220 2748 9222
rect 2804 9220 2828 9222
rect 2884 9220 2890 9222
rect 2582 9200 2890 9220
rect 2582 8188 2890 8208
rect 2582 8186 2588 8188
rect 2644 8186 2668 8188
rect 2724 8186 2748 8188
rect 2804 8186 2828 8188
rect 2884 8186 2890 8188
rect 2644 8134 2646 8186
rect 2826 8134 2828 8186
rect 2582 8132 2588 8134
rect 2644 8132 2668 8134
rect 2724 8132 2748 8134
rect 2804 8132 2828 8134
rect 2884 8132 2890 8134
rect 2582 8112 2890 8132
rect 2582 7100 2890 7120
rect 2582 7098 2588 7100
rect 2644 7098 2668 7100
rect 2724 7098 2748 7100
rect 2804 7098 2828 7100
rect 2884 7098 2890 7100
rect 2644 7046 2646 7098
rect 2826 7046 2828 7098
rect 2582 7044 2588 7046
rect 2644 7044 2668 7046
rect 2724 7044 2748 7046
rect 2804 7044 2828 7046
rect 2884 7044 2890 7046
rect 2582 7024 2890 7044
rect 2976 6798 3004 11018
rect 3252 10810 3280 24754
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3608 23520 3660 23526
rect 3608 23462 3660 23468
rect 3424 23044 3476 23050
rect 3424 22986 3476 22992
rect 3330 22128 3386 22137
rect 3330 22063 3386 22072
rect 3344 21554 3372 22063
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3344 18290 3372 20198
rect 3436 19242 3464 22986
rect 3620 22098 3648 23462
rect 3804 22681 3832 23666
rect 3896 22778 3924 24346
rect 3884 22772 3936 22778
rect 3884 22714 3936 22720
rect 3790 22672 3846 22681
rect 3790 22607 3846 22616
rect 3608 22092 3660 22098
rect 3608 22034 3660 22040
rect 3792 21344 3844 21350
rect 3792 21286 3844 21292
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3528 20369 3556 20402
rect 3514 20360 3570 20369
rect 3514 20295 3570 20304
rect 3516 19916 3568 19922
rect 3516 19858 3568 19864
rect 3424 19236 3476 19242
rect 3424 19178 3476 19184
rect 3528 18970 3556 19858
rect 3804 19854 3832 21286
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 3988 19514 4016 26206
rect 4213 26140 4521 26160
rect 4213 26138 4219 26140
rect 4275 26138 4299 26140
rect 4355 26138 4379 26140
rect 4435 26138 4459 26140
rect 4515 26138 4521 26140
rect 4275 26086 4277 26138
rect 4457 26086 4459 26138
rect 4213 26084 4219 26086
rect 4275 26084 4299 26086
rect 4355 26084 4379 26086
rect 4435 26084 4459 26086
rect 4515 26084 4521 26086
rect 4213 26064 4521 26084
rect 4068 25356 4120 25362
rect 4068 25298 4120 25304
rect 4080 23866 4108 25298
rect 4213 25052 4521 25072
rect 4213 25050 4219 25052
rect 4275 25050 4299 25052
rect 4355 25050 4379 25052
rect 4435 25050 4459 25052
rect 4515 25050 4521 25052
rect 4275 24998 4277 25050
rect 4457 24998 4459 25050
rect 4213 24996 4219 24998
rect 4275 24996 4299 24998
rect 4355 24996 4379 24998
rect 4435 24996 4459 24998
rect 4515 24996 4521 24998
rect 4213 24976 4521 24996
rect 4252 24812 4304 24818
rect 4252 24754 4304 24760
rect 4264 24206 4292 24754
rect 4632 24342 4660 27798
rect 4724 24410 4752 55558
rect 4802 51640 4858 51649
rect 4802 51575 4858 51584
rect 4816 40730 4844 51575
rect 4908 51074 4936 61134
rect 5000 51241 5028 73510
rect 5080 65136 5132 65142
rect 5080 65078 5132 65084
rect 4986 51232 5042 51241
rect 4986 51167 5042 51176
rect 4908 51046 5028 51074
rect 4894 50960 4950 50969
rect 4894 50895 4950 50904
rect 4908 47190 4936 50895
rect 4896 47184 4948 47190
rect 4896 47126 4948 47132
rect 4896 46368 4948 46374
rect 4896 46310 4948 46316
rect 4908 42294 4936 46310
rect 5000 43382 5028 51046
rect 5092 46170 5120 65078
rect 5184 52630 5212 74802
rect 5845 74556 6153 74576
rect 5845 74554 5851 74556
rect 5907 74554 5931 74556
rect 5987 74554 6011 74556
rect 6067 74554 6091 74556
rect 6147 74554 6153 74556
rect 5907 74502 5909 74554
rect 6089 74502 6091 74554
rect 5845 74500 5851 74502
rect 5907 74500 5931 74502
rect 5987 74500 6011 74502
rect 6067 74500 6091 74502
rect 6147 74500 6153 74502
rect 5845 74480 6153 74500
rect 9109 74556 9417 74576
rect 9109 74554 9115 74556
rect 9171 74554 9195 74556
rect 9251 74554 9275 74556
rect 9331 74554 9355 74556
rect 9411 74554 9417 74556
rect 9171 74502 9173 74554
rect 9353 74502 9355 74554
rect 9109 74500 9115 74502
rect 9171 74500 9195 74502
rect 9251 74500 9275 74502
rect 9331 74500 9355 74502
rect 9411 74500 9417 74502
rect 9109 74480 9417 74500
rect 8300 74384 8352 74390
rect 8300 74326 8352 74332
rect 7477 74012 7785 74032
rect 7477 74010 7483 74012
rect 7539 74010 7563 74012
rect 7619 74010 7643 74012
rect 7699 74010 7723 74012
rect 7779 74010 7785 74012
rect 7539 73958 7541 74010
rect 7721 73958 7723 74010
rect 7477 73956 7483 73958
rect 7539 73956 7563 73958
rect 7619 73956 7643 73958
rect 7699 73956 7723 73958
rect 7779 73956 7785 73958
rect 7477 73936 7785 73956
rect 5845 73468 6153 73488
rect 5845 73466 5851 73468
rect 5907 73466 5931 73468
rect 5987 73466 6011 73468
rect 6067 73466 6091 73468
rect 6147 73466 6153 73468
rect 5907 73414 5909 73466
rect 6089 73414 6091 73466
rect 5845 73412 5851 73414
rect 5907 73412 5931 73414
rect 5987 73412 6011 73414
rect 6067 73412 6091 73414
rect 6147 73412 6153 73414
rect 5845 73392 6153 73412
rect 5540 73160 5592 73166
rect 5540 73102 5592 73108
rect 5264 70440 5316 70446
rect 5264 70382 5316 70388
rect 5276 53242 5304 70382
rect 5356 59628 5408 59634
rect 5356 59570 5408 59576
rect 5264 53236 5316 53242
rect 5264 53178 5316 53184
rect 5368 53145 5396 59570
rect 5448 59016 5500 59022
rect 5448 58958 5500 58964
rect 5460 53689 5488 58958
rect 5446 53680 5502 53689
rect 5446 53615 5502 53624
rect 5448 53576 5500 53582
rect 5448 53518 5500 53524
rect 5354 53136 5410 53145
rect 5264 53100 5316 53106
rect 5354 53071 5410 53080
rect 5264 53042 5316 53048
rect 5172 52624 5224 52630
rect 5172 52566 5224 52572
rect 5276 51898 5304 53042
rect 5356 52964 5408 52970
rect 5356 52906 5408 52912
rect 5184 51870 5304 51898
rect 5184 51082 5212 51870
rect 5368 51377 5396 52906
rect 5354 51368 5410 51377
rect 5354 51303 5410 51312
rect 5460 51218 5488 53518
rect 5552 51542 5580 73102
rect 7477 72924 7785 72944
rect 7477 72922 7483 72924
rect 7539 72922 7563 72924
rect 7619 72922 7643 72924
rect 7699 72922 7723 72924
rect 7779 72922 7785 72924
rect 7539 72870 7541 72922
rect 7721 72870 7723 72922
rect 7477 72868 7483 72870
rect 7539 72868 7563 72870
rect 7619 72868 7643 72870
rect 7699 72868 7723 72870
rect 7779 72868 7785 72870
rect 7477 72848 7785 72868
rect 5845 72380 6153 72400
rect 5845 72378 5851 72380
rect 5907 72378 5931 72380
rect 5987 72378 6011 72380
rect 6067 72378 6091 72380
rect 6147 72378 6153 72380
rect 5907 72326 5909 72378
rect 6089 72326 6091 72378
rect 5845 72324 5851 72326
rect 5907 72324 5931 72326
rect 5987 72324 6011 72326
rect 6067 72324 6091 72326
rect 6147 72324 6153 72326
rect 5845 72304 6153 72324
rect 7477 71836 7785 71856
rect 7477 71834 7483 71836
rect 7539 71834 7563 71836
rect 7619 71834 7643 71836
rect 7699 71834 7723 71836
rect 7779 71834 7785 71836
rect 7539 71782 7541 71834
rect 7721 71782 7723 71834
rect 7477 71780 7483 71782
rect 7539 71780 7563 71782
rect 7619 71780 7643 71782
rect 7699 71780 7723 71782
rect 7779 71780 7785 71782
rect 7477 71760 7785 71780
rect 5845 71292 6153 71312
rect 5845 71290 5851 71292
rect 5907 71290 5931 71292
rect 5987 71290 6011 71292
rect 6067 71290 6091 71292
rect 6147 71290 6153 71292
rect 5907 71238 5909 71290
rect 6089 71238 6091 71290
rect 5845 71236 5851 71238
rect 5907 71236 5931 71238
rect 5987 71236 6011 71238
rect 6067 71236 6091 71238
rect 6147 71236 6153 71238
rect 5845 71216 6153 71236
rect 7477 70748 7785 70768
rect 7477 70746 7483 70748
rect 7539 70746 7563 70748
rect 7619 70746 7643 70748
rect 7699 70746 7723 70748
rect 7779 70746 7785 70748
rect 7539 70694 7541 70746
rect 7721 70694 7723 70746
rect 7477 70692 7483 70694
rect 7539 70692 7563 70694
rect 7619 70692 7643 70694
rect 7699 70692 7723 70694
rect 7779 70692 7785 70694
rect 7477 70672 7785 70692
rect 5845 70204 6153 70224
rect 5845 70202 5851 70204
rect 5907 70202 5931 70204
rect 5987 70202 6011 70204
rect 6067 70202 6091 70204
rect 6147 70202 6153 70204
rect 5907 70150 5909 70202
rect 6089 70150 6091 70202
rect 5845 70148 5851 70150
rect 5907 70148 5931 70150
rect 5987 70148 6011 70150
rect 6067 70148 6091 70150
rect 6147 70148 6153 70150
rect 5845 70128 6153 70148
rect 7477 69660 7785 69680
rect 7477 69658 7483 69660
rect 7539 69658 7563 69660
rect 7619 69658 7643 69660
rect 7699 69658 7723 69660
rect 7779 69658 7785 69660
rect 7539 69606 7541 69658
rect 7721 69606 7723 69658
rect 7477 69604 7483 69606
rect 7539 69604 7563 69606
rect 7619 69604 7643 69606
rect 7699 69604 7723 69606
rect 7779 69604 7785 69606
rect 7477 69584 7785 69604
rect 5845 69116 6153 69136
rect 5845 69114 5851 69116
rect 5907 69114 5931 69116
rect 5987 69114 6011 69116
rect 6067 69114 6091 69116
rect 6147 69114 6153 69116
rect 5907 69062 5909 69114
rect 6089 69062 6091 69114
rect 5845 69060 5851 69062
rect 5907 69060 5931 69062
rect 5987 69060 6011 69062
rect 6067 69060 6091 69062
rect 6147 69060 6153 69062
rect 5845 69040 6153 69060
rect 7477 68572 7785 68592
rect 7477 68570 7483 68572
rect 7539 68570 7563 68572
rect 7619 68570 7643 68572
rect 7699 68570 7723 68572
rect 7779 68570 7785 68572
rect 7539 68518 7541 68570
rect 7721 68518 7723 68570
rect 7477 68516 7483 68518
rect 7539 68516 7563 68518
rect 7619 68516 7643 68518
rect 7699 68516 7723 68518
rect 7779 68516 7785 68518
rect 7477 68496 7785 68516
rect 5845 68028 6153 68048
rect 5845 68026 5851 68028
rect 5907 68026 5931 68028
rect 5987 68026 6011 68028
rect 6067 68026 6091 68028
rect 6147 68026 6153 68028
rect 5907 67974 5909 68026
rect 6089 67974 6091 68026
rect 5845 67972 5851 67974
rect 5907 67972 5931 67974
rect 5987 67972 6011 67974
rect 6067 67972 6091 67974
rect 6147 67972 6153 67974
rect 5845 67952 6153 67972
rect 6920 67856 6972 67862
rect 6920 67798 6972 67804
rect 5845 66940 6153 66960
rect 5845 66938 5851 66940
rect 5907 66938 5931 66940
rect 5987 66938 6011 66940
rect 6067 66938 6091 66940
rect 6147 66938 6153 66940
rect 5907 66886 5909 66938
rect 6089 66886 6091 66938
rect 5845 66884 5851 66886
rect 5907 66884 5931 66886
rect 5987 66884 6011 66886
rect 6067 66884 6091 66886
rect 6147 66884 6153 66886
rect 5845 66864 6153 66884
rect 5845 65852 6153 65872
rect 5845 65850 5851 65852
rect 5907 65850 5931 65852
rect 5987 65850 6011 65852
rect 6067 65850 6091 65852
rect 6147 65850 6153 65852
rect 5907 65798 5909 65850
rect 6089 65798 6091 65850
rect 5845 65796 5851 65798
rect 5907 65796 5931 65798
rect 5987 65796 6011 65798
rect 6067 65796 6091 65798
rect 6147 65796 6153 65798
rect 5845 65776 6153 65796
rect 5845 64764 6153 64784
rect 5845 64762 5851 64764
rect 5907 64762 5931 64764
rect 5987 64762 6011 64764
rect 6067 64762 6091 64764
rect 6147 64762 6153 64764
rect 5907 64710 5909 64762
rect 6089 64710 6091 64762
rect 5845 64708 5851 64710
rect 5907 64708 5931 64710
rect 5987 64708 6011 64710
rect 6067 64708 6091 64710
rect 6147 64708 6153 64710
rect 5845 64688 6153 64708
rect 6736 63776 6788 63782
rect 6736 63718 6788 63724
rect 5845 63676 6153 63696
rect 5845 63674 5851 63676
rect 5907 63674 5931 63676
rect 5987 63674 6011 63676
rect 6067 63674 6091 63676
rect 6147 63674 6153 63676
rect 5907 63622 5909 63674
rect 6089 63622 6091 63674
rect 5845 63620 5851 63622
rect 5907 63620 5931 63622
rect 5987 63620 6011 63622
rect 6067 63620 6091 63622
rect 6147 63620 6153 63622
rect 5845 63600 6153 63620
rect 5724 63368 5776 63374
rect 5724 63310 5776 63316
rect 5632 61124 5684 61130
rect 5632 61066 5684 61072
rect 5540 51536 5592 51542
rect 5540 51478 5592 51484
rect 5460 51190 5580 51218
rect 5446 51096 5502 51105
rect 5184 51054 5304 51082
rect 5172 50924 5224 50930
rect 5172 50866 5224 50872
rect 5080 46164 5132 46170
rect 5080 46106 5132 46112
rect 4988 43376 5040 43382
rect 4988 43318 5040 43324
rect 4988 42696 5040 42702
rect 4988 42638 5040 42644
rect 4896 42288 4948 42294
rect 4896 42230 4948 42236
rect 5000 42226 5028 42638
rect 5080 42288 5132 42294
rect 5080 42230 5132 42236
rect 4988 42220 5040 42226
rect 4988 42162 5040 42168
rect 4896 41200 4948 41206
rect 4896 41142 4948 41148
rect 4804 40724 4856 40730
rect 4804 40666 4856 40672
rect 4804 40112 4856 40118
rect 4804 40054 4856 40060
rect 4816 38894 4844 40054
rect 4804 38888 4856 38894
rect 4804 38830 4856 38836
rect 4816 36922 4844 38830
rect 4804 36916 4856 36922
rect 4804 36858 4856 36864
rect 4804 35080 4856 35086
rect 4804 35022 4856 35028
rect 4816 32366 4844 35022
rect 4908 33386 4936 41142
rect 5000 41138 5028 42162
rect 4988 41132 5040 41138
rect 4988 41074 5040 41080
rect 4896 33380 4948 33386
rect 4896 33322 4948 33328
rect 4896 32836 4948 32842
rect 4896 32778 4948 32784
rect 4804 32360 4856 32366
rect 4804 32302 4856 32308
rect 4816 28082 4844 32302
rect 4908 30666 4936 32778
rect 4896 30660 4948 30666
rect 4896 30602 4948 30608
rect 4908 29714 4936 30602
rect 4896 29708 4948 29714
rect 4896 29650 4948 29656
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 5000 24614 5028 41074
rect 5092 34746 5120 42230
rect 5080 34740 5132 34746
rect 5080 34682 5132 34688
rect 4988 24608 5040 24614
rect 4988 24550 5040 24556
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 4620 24336 4672 24342
rect 4620 24278 4672 24284
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 4213 23964 4521 23984
rect 4213 23962 4219 23964
rect 4275 23962 4299 23964
rect 4355 23962 4379 23964
rect 4435 23962 4459 23964
rect 4515 23962 4521 23964
rect 4275 23910 4277 23962
rect 4457 23910 4459 23962
rect 4213 23908 4219 23910
rect 4275 23908 4299 23910
rect 4355 23908 4379 23910
rect 4435 23908 4459 23910
rect 4515 23908 4521 23910
rect 4213 23888 4521 23908
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4344 23792 4396 23798
rect 4344 23734 4396 23740
rect 4068 23656 4120 23662
rect 4068 23598 4120 23604
rect 4080 23118 4108 23598
rect 4356 23118 4384 23734
rect 4632 23338 4660 24278
rect 4632 23310 4844 23338
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4213 22876 4521 22896
rect 4213 22874 4219 22876
rect 4275 22874 4299 22876
rect 4355 22874 4379 22876
rect 4435 22874 4459 22876
rect 4515 22874 4521 22876
rect 4275 22822 4277 22874
rect 4457 22822 4459 22874
rect 4213 22820 4219 22822
rect 4275 22820 4299 22822
rect 4355 22820 4379 22822
rect 4435 22820 4459 22822
rect 4515 22820 4521 22822
rect 4213 22800 4521 22820
rect 4632 22642 4660 23122
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4724 22778 4752 22918
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4632 22030 4660 22578
rect 4816 22574 4844 23310
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 4712 22500 4764 22506
rect 4712 22442 4764 22448
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4213 21788 4521 21808
rect 4213 21786 4219 21788
rect 4275 21786 4299 21788
rect 4355 21786 4379 21788
rect 4435 21786 4459 21788
rect 4515 21786 4521 21788
rect 4275 21734 4277 21786
rect 4457 21734 4459 21786
rect 4213 21732 4219 21734
rect 4275 21732 4299 21734
rect 4355 21732 4379 21734
rect 4435 21732 4459 21734
rect 4515 21732 4521 21734
rect 4213 21712 4521 21732
rect 4632 21554 4660 21966
rect 4724 21554 4752 22442
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4816 21010 4844 22510
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4908 21146 4936 21286
rect 4896 21140 4948 21146
rect 4896 21082 4948 21088
rect 5000 21026 5028 24550
rect 4804 21004 4856 21010
rect 4804 20946 4856 20952
rect 4908 20998 5028 21026
rect 4712 20936 4764 20942
rect 4712 20878 4764 20884
rect 4213 20700 4521 20720
rect 4213 20698 4219 20700
rect 4275 20698 4299 20700
rect 4355 20698 4379 20700
rect 4435 20698 4459 20700
rect 4515 20698 4521 20700
rect 4275 20646 4277 20698
rect 4457 20646 4459 20698
rect 4213 20644 4219 20646
rect 4275 20644 4299 20646
rect 4355 20644 4379 20646
rect 4435 20644 4459 20646
rect 4515 20644 4521 20646
rect 4213 20624 4521 20644
rect 4160 20528 4212 20534
rect 4160 20470 4212 20476
rect 4172 19802 4200 20470
rect 4620 20324 4672 20330
rect 4620 20266 4672 20272
rect 4080 19774 4200 19802
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4080 19378 4108 19774
rect 4213 19612 4521 19632
rect 4213 19610 4219 19612
rect 4275 19610 4299 19612
rect 4355 19610 4379 19612
rect 4435 19610 4459 19612
rect 4515 19610 4521 19612
rect 4275 19558 4277 19610
rect 4457 19558 4459 19610
rect 4213 19556 4219 19558
rect 4275 19556 4299 19558
rect 4355 19556 4379 19558
rect 4435 19556 4459 19558
rect 4515 19556 4521 19558
rect 4213 19536 4521 19556
rect 4632 19446 4660 20266
rect 4620 19440 4672 19446
rect 4620 19382 4672 19388
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3528 18850 3556 18906
rect 3436 18822 3556 18850
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3344 16590 3372 18022
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3436 11762 3464 18822
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3792 18624 3844 18630
rect 3988 18601 4016 18702
rect 3792 18566 3844 18572
rect 3974 18592 4030 18601
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3528 18193 3556 18226
rect 3514 18184 3570 18193
rect 3514 18119 3570 18128
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3712 9586 3740 17274
rect 3804 17202 3832 18566
rect 3974 18527 4030 18536
rect 4213 18524 4521 18544
rect 4213 18522 4219 18524
rect 4275 18522 4299 18524
rect 4355 18522 4379 18524
rect 4435 18522 4459 18524
rect 4515 18522 4521 18524
rect 4275 18470 4277 18522
rect 4457 18470 4459 18522
rect 4213 18468 4219 18470
rect 4275 18468 4299 18470
rect 4355 18468 4379 18470
rect 4435 18468 4459 18470
rect 4515 18468 4521 18470
rect 4213 18448 4521 18468
rect 4632 18358 4660 19382
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 4724 18290 4752 20878
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4712 18284 4764 18290
rect 4712 18226 4764 18232
rect 4344 18148 4396 18154
rect 4344 18090 4396 18096
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3896 7886 3924 11154
rect 3988 10062 4016 17818
rect 4356 17678 4384 18090
rect 4724 17678 4752 18226
rect 4344 17672 4396 17678
rect 4344 17614 4396 17620
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4213 17436 4521 17456
rect 4213 17434 4219 17436
rect 4275 17434 4299 17436
rect 4355 17434 4379 17436
rect 4435 17434 4459 17436
rect 4515 17434 4521 17436
rect 4275 17382 4277 17434
rect 4457 17382 4459 17434
rect 4213 17380 4219 17382
rect 4275 17380 4299 17382
rect 4355 17380 4379 17382
rect 4435 17380 4459 17382
rect 4515 17380 4521 17382
rect 4213 17360 4521 17380
rect 4724 17202 4752 17614
rect 4816 17270 4844 19314
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4213 16348 4521 16368
rect 4213 16346 4219 16348
rect 4275 16346 4299 16348
rect 4355 16346 4379 16348
rect 4435 16346 4459 16348
rect 4515 16346 4521 16348
rect 4275 16294 4277 16346
rect 4457 16294 4459 16346
rect 4213 16292 4219 16294
rect 4275 16292 4299 16294
rect 4355 16292 4379 16294
rect 4435 16292 4459 16294
rect 4515 16292 4521 16294
rect 4213 16272 4521 16292
rect 4213 15260 4521 15280
rect 4213 15258 4219 15260
rect 4275 15258 4299 15260
rect 4355 15258 4379 15260
rect 4435 15258 4459 15260
rect 4515 15258 4521 15260
rect 4275 15206 4277 15258
rect 4457 15206 4459 15258
rect 4213 15204 4219 15206
rect 4275 15204 4299 15206
rect 4355 15204 4379 15206
rect 4435 15204 4459 15206
rect 4515 15204 4521 15206
rect 4213 15184 4521 15204
rect 4213 14172 4521 14192
rect 4213 14170 4219 14172
rect 4275 14170 4299 14172
rect 4355 14170 4379 14172
rect 4435 14170 4459 14172
rect 4515 14170 4521 14172
rect 4275 14118 4277 14170
rect 4457 14118 4459 14170
rect 4213 14116 4219 14118
rect 4275 14116 4299 14118
rect 4355 14116 4379 14118
rect 4435 14116 4459 14118
rect 4515 14116 4521 14118
rect 4213 14096 4521 14116
rect 4213 13084 4521 13104
rect 4213 13082 4219 13084
rect 4275 13082 4299 13084
rect 4355 13082 4379 13084
rect 4435 13082 4459 13084
rect 4515 13082 4521 13084
rect 4275 13030 4277 13082
rect 4457 13030 4459 13082
rect 4213 13028 4219 13030
rect 4275 13028 4299 13030
rect 4355 13028 4379 13030
rect 4435 13028 4459 13030
rect 4515 13028 4521 13030
rect 4213 13008 4521 13028
rect 4213 11996 4521 12016
rect 4213 11994 4219 11996
rect 4275 11994 4299 11996
rect 4355 11994 4379 11996
rect 4435 11994 4459 11996
rect 4515 11994 4521 11996
rect 4275 11942 4277 11994
rect 4457 11942 4459 11994
rect 4213 11940 4219 11942
rect 4275 11940 4299 11942
rect 4355 11940 4379 11942
rect 4435 11940 4459 11942
rect 4515 11940 4521 11942
rect 4213 11920 4521 11940
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4172 11150 4200 11698
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4213 10908 4521 10928
rect 4213 10906 4219 10908
rect 4275 10906 4299 10908
rect 4355 10906 4379 10908
rect 4435 10906 4459 10908
rect 4515 10906 4521 10908
rect 4275 10854 4277 10906
rect 4457 10854 4459 10906
rect 4213 10852 4219 10854
rect 4275 10852 4299 10854
rect 4355 10852 4379 10854
rect 4435 10852 4459 10854
rect 4515 10852 4521 10854
rect 4213 10832 4521 10852
rect 4632 10606 4660 11086
rect 4908 10674 4936 20998
rect 5184 19922 5212 50866
rect 5276 41546 5304 51054
rect 5446 51031 5502 51040
rect 5354 50960 5410 50969
rect 5354 50895 5410 50904
rect 5264 41540 5316 41546
rect 5264 41482 5316 41488
rect 5262 41440 5318 41449
rect 5262 41375 5318 41384
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 4988 19780 5040 19786
rect 4988 19722 5040 19728
rect 5000 17678 5028 19722
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5000 17338 5028 17478
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 5276 11218 5304 41375
rect 5368 41206 5396 50895
rect 5460 50810 5488 51031
rect 5552 50930 5580 51190
rect 5540 50924 5592 50930
rect 5540 50866 5592 50872
rect 5460 50782 5580 50810
rect 5448 50720 5500 50726
rect 5448 50662 5500 50668
rect 5460 42634 5488 50662
rect 5552 45558 5580 50782
rect 5540 45552 5592 45558
rect 5540 45494 5592 45500
rect 5448 42628 5500 42634
rect 5448 42570 5500 42576
rect 5356 41200 5408 41206
rect 5356 41142 5408 41148
rect 5356 40724 5408 40730
rect 5356 40666 5408 40672
rect 5368 33046 5396 40666
rect 5460 34678 5488 42570
rect 5448 34672 5500 34678
rect 5448 34614 5500 34620
rect 5644 33862 5672 61066
rect 5736 39574 5764 63310
rect 5845 62588 6153 62608
rect 5845 62586 5851 62588
rect 5907 62586 5931 62588
rect 5987 62586 6011 62588
rect 6067 62586 6091 62588
rect 6147 62586 6153 62588
rect 5907 62534 5909 62586
rect 6089 62534 6091 62586
rect 5845 62532 5851 62534
rect 5907 62532 5931 62534
rect 5987 62532 6011 62534
rect 6067 62532 6091 62534
rect 6147 62532 6153 62534
rect 5845 62512 6153 62532
rect 5845 61500 6153 61520
rect 5845 61498 5851 61500
rect 5907 61498 5931 61500
rect 5987 61498 6011 61500
rect 6067 61498 6091 61500
rect 6147 61498 6153 61500
rect 5907 61446 5909 61498
rect 6089 61446 6091 61498
rect 5845 61444 5851 61446
rect 5907 61444 5931 61446
rect 5987 61444 6011 61446
rect 6067 61444 6091 61446
rect 6147 61444 6153 61446
rect 5845 61424 6153 61444
rect 5845 60412 6153 60432
rect 5845 60410 5851 60412
rect 5907 60410 5931 60412
rect 5987 60410 6011 60412
rect 6067 60410 6091 60412
rect 6147 60410 6153 60412
rect 5907 60358 5909 60410
rect 6089 60358 6091 60410
rect 5845 60356 5851 60358
rect 5907 60356 5931 60358
rect 5987 60356 6011 60358
rect 6067 60356 6091 60358
rect 6147 60356 6153 60358
rect 5845 60336 6153 60356
rect 6276 60104 6328 60110
rect 6276 60046 6328 60052
rect 5845 59324 6153 59344
rect 5845 59322 5851 59324
rect 5907 59322 5931 59324
rect 5987 59322 6011 59324
rect 6067 59322 6091 59324
rect 6147 59322 6153 59324
rect 5907 59270 5909 59322
rect 6089 59270 6091 59322
rect 5845 59268 5851 59270
rect 5907 59268 5931 59270
rect 5987 59268 6011 59270
rect 6067 59268 6091 59270
rect 6147 59268 6153 59270
rect 5845 59248 6153 59268
rect 5845 58236 6153 58256
rect 5845 58234 5851 58236
rect 5907 58234 5931 58236
rect 5987 58234 6011 58236
rect 6067 58234 6091 58236
rect 6147 58234 6153 58236
rect 5907 58182 5909 58234
rect 6089 58182 6091 58234
rect 5845 58180 5851 58182
rect 5907 58180 5931 58182
rect 5987 58180 6011 58182
rect 6067 58180 6091 58182
rect 6147 58180 6153 58182
rect 5845 58160 6153 58180
rect 6184 57452 6236 57458
rect 6184 57394 6236 57400
rect 5845 57148 6153 57168
rect 5845 57146 5851 57148
rect 5907 57146 5931 57148
rect 5987 57146 6011 57148
rect 6067 57146 6091 57148
rect 6147 57146 6153 57148
rect 5907 57094 5909 57146
rect 6089 57094 6091 57146
rect 5845 57092 5851 57094
rect 5907 57092 5931 57094
rect 5987 57092 6011 57094
rect 6067 57092 6091 57094
rect 6147 57092 6153 57094
rect 5845 57072 6153 57092
rect 5845 56060 6153 56080
rect 5845 56058 5851 56060
rect 5907 56058 5931 56060
rect 5987 56058 6011 56060
rect 6067 56058 6091 56060
rect 6147 56058 6153 56060
rect 5907 56006 5909 56058
rect 6089 56006 6091 56058
rect 5845 56004 5851 56006
rect 5907 56004 5931 56006
rect 5987 56004 6011 56006
rect 6067 56004 6091 56006
rect 6147 56004 6153 56006
rect 5845 55984 6153 56004
rect 5845 54972 6153 54992
rect 5845 54970 5851 54972
rect 5907 54970 5931 54972
rect 5987 54970 6011 54972
rect 6067 54970 6091 54972
rect 6147 54970 6153 54972
rect 5907 54918 5909 54970
rect 6089 54918 6091 54970
rect 5845 54916 5851 54918
rect 5907 54916 5931 54918
rect 5987 54916 6011 54918
rect 6067 54916 6091 54918
rect 6147 54916 6153 54918
rect 5845 54896 6153 54916
rect 5845 53884 6153 53904
rect 5845 53882 5851 53884
rect 5907 53882 5931 53884
rect 5987 53882 6011 53884
rect 6067 53882 6091 53884
rect 6147 53882 6153 53884
rect 5907 53830 5909 53882
rect 6089 53830 6091 53882
rect 5845 53828 5851 53830
rect 5907 53828 5931 53830
rect 5987 53828 6011 53830
rect 6067 53828 6091 53830
rect 6147 53828 6153 53830
rect 5845 53808 6153 53828
rect 5845 52796 6153 52816
rect 5845 52794 5851 52796
rect 5907 52794 5931 52796
rect 5987 52794 6011 52796
rect 6067 52794 6091 52796
rect 6147 52794 6153 52796
rect 5907 52742 5909 52794
rect 6089 52742 6091 52794
rect 5845 52740 5851 52742
rect 5907 52740 5931 52742
rect 5987 52740 6011 52742
rect 6067 52740 6091 52742
rect 6147 52740 6153 52742
rect 5845 52720 6153 52740
rect 5845 51708 6153 51728
rect 5845 51706 5851 51708
rect 5907 51706 5931 51708
rect 5987 51706 6011 51708
rect 6067 51706 6091 51708
rect 6147 51706 6153 51708
rect 5907 51654 5909 51706
rect 6089 51654 6091 51706
rect 5845 51652 5851 51654
rect 5907 51652 5931 51654
rect 5987 51652 6011 51654
rect 6067 51652 6091 51654
rect 6147 51652 6153 51654
rect 5845 51632 6153 51652
rect 5816 51536 5868 51542
rect 5816 51478 5868 51484
rect 5828 50794 5856 51478
rect 5816 50788 5868 50794
rect 5816 50730 5868 50736
rect 5845 50620 6153 50640
rect 5845 50618 5851 50620
rect 5907 50618 5931 50620
rect 5987 50618 6011 50620
rect 6067 50618 6091 50620
rect 6147 50618 6153 50620
rect 5907 50566 5909 50618
rect 6089 50566 6091 50618
rect 5845 50564 5851 50566
rect 5907 50564 5931 50566
rect 5987 50564 6011 50566
rect 6067 50564 6091 50566
rect 6147 50564 6153 50566
rect 5845 50544 6153 50564
rect 5845 49532 6153 49552
rect 5845 49530 5851 49532
rect 5907 49530 5931 49532
rect 5987 49530 6011 49532
rect 6067 49530 6091 49532
rect 6147 49530 6153 49532
rect 5907 49478 5909 49530
rect 6089 49478 6091 49530
rect 5845 49476 5851 49478
rect 5907 49476 5931 49478
rect 5987 49476 6011 49478
rect 6067 49476 6091 49478
rect 6147 49476 6153 49478
rect 5845 49456 6153 49476
rect 5845 48444 6153 48464
rect 5845 48442 5851 48444
rect 5907 48442 5931 48444
rect 5987 48442 6011 48444
rect 6067 48442 6091 48444
rect 6147 48442 6153 48444
rect 5907 48390 5909 48442
rect 6089 48390 6091 48442
rect 5845 48388 5851 48390
rect 5907 48388 5931 48390
rect 5987 48388 6011 48390
rect 6067 48388 6091 48390
rect 6147 48388 6153 48390
rect 5845 48368 6153 48388
rect 5845 47356 6153 47376
rect 5845 47354 5851 47356
rect 5907 47354 5931 47356
rect 5987 47354 6011 47356
rect 6067 47354 6091 47356
rect 6147 47354 6153 47356
rect 5907 47302 5909 47354
rect 6089 47302 6091 47354
rect 5845 47300 5851 47302
rect 5907 47300 5931 47302
rect 5987 47300 6011 47302
rect 6067 47300 6091 47302
rect 6147 47300 6153 47302
rect 5845 47280 6153 47300
rect 5845 46268 6153 46288
rect 5845 46266 5851 46268
rect 5907 46266 5931 46268
rect 5987 46266 6011 46268
rect 6067 46266 6091 46268
rect 6147 46266 6153 46268
rect 5907 46214 5909 46266
rect 6089 46214 6091 46266
rect 5845 46212 5851 46214
rect 5907 46212 5931 46214
rect 5987 46212 6011 46214
rect 6067 46212 6091 46214
rect 6147 46212 6153 46214
rect 5845 46192 6153 46212
rect 5845 45180 6153 45200
rect 5845 45178 5851 45180
rect 5907 45178 5931 45180
rect 5987 45178 6011 45180
rect 6067 45178 6091 45180
rect 6147 45178 6153 45180
rect 5907 45126 5909 45178
rect 6089 45126 6091 45178
rect 5845 45124 5851 45126
rect 5907 45124 5931 45126
rect 5987 45124 6011 45126
rect 6067 45124 6091 45126
rect 6147 45124 6153 45126
rect 5845 45104 6153 45124
rect 5845 44092 6153 44112
rect 5845 44090 5851 44092
rect 5907 44090 5931 44092
rect 5987 44090 6011 44092
rect 6067 44090 6091 44092
rect 6147 44090 6153 44092
rect 5907 44038 5909 44090
rect 6089 44038 6091 44090
rect 5845 44036 5851 44038
rect 5907 44036 5931 44038
rect 5987 44036 6011 44038
rect 6067 44036 6091 44038
rect 6147 44036 6153 44038
rect 5845 44016 6153 44036
rect 5845 43004 6153 43024
rect 5845 43002 5851 43004
rect 5907 43002 5931 43004
rect 5987 43002 6011 43004
rect 6067 43002 6091 43004
rect 6147 43002 6153 43004
rect 5907 42950 5909 43002
rect 6089 42950 6091 43002
rect 5845 42948 5851 42950
rect 5907 42948 5931 42950
rect 5987 42948 6011 42950
rect 6067 42948 6091 42950
rect 6147 42948 6153 42950
rect 5845 42928 6153 42948
rect 5845 41916 6153 41936
rect 5845 41914 5851 41916
rect 5907 41914 5931 41916
rect 5987 41914 6011 41916
rect 6067 41914 6091 41916
rect 6147 41914 6153 41916
rect 5907 41862 5909 41914
rect 6089 41862 6091 41914
rect 5845 41860 5851 41862
rect 5907 41860 5931 41862
rect 5987 41860 6011 41862
rect 6067 41860 6091 41862
rect 6147 41860 6153 41862
rect 5845 41840 6153 41860
rect 5845 40828 6153 40848
rect 5845 40826 5851 40828
rect 5907 40826 5931 40828
rect 5987 40826 6011 40828
rect 6067 40826 6091 40828
rect 6147 40826 6153 40828
rect 5907 40774 5909 40826
rect 6089 40774 6091 40826
rect 5845 40772 5851 40774
rect 5907 40772 5931 40774
rect 5987 40772 6011 40774
rect 6067 40772 6091 40774
rect 6147 40772 6153 40774
rect 5845 40752 6153 40772
rect 5845 39740 6153 39760
rect 5845 39738 5851 39740
rect 5907 39738 5931 39740
rect 5987 39738 6011 39740
rect 6067 39738 6091 39740
rect 6147 39738 6153 39740
rect 5907 39686 5909 39738
rect 6089 39686 6091 39738
rect 5845 39684 5851 39686
rect 5907 39684 5931 39686
rect 5987 39684 6011 39686
rect 6067 39684 6091 39686
rect 6147 39684 6153 39686
rect 5845 39664 6153 39684
rect 5724 39568 5776 39574
rect 5724 39510 5776 39516
rect 5845 38652 6153 38672
rect 5845 38650 5851 38652
rect 5907 38650 5931 38652
rect 5987 38650 6011 38652
rect 6067 38650 6091 38652
rect 6147 38650 6153 38652
rect 5907 38598 5909 38650
rect 6089 38598 6091 38650
rect 5845 38596 5851 38598
rect 5907 38596 5931 38598
rect 5987 38596 6011 38598
rect 6067 38596 6091 38598
rect 6147 38596 6153 38598
rect 5845 38576 6153 38596
rect 5845 37564 6153 37584
rect 5845 37562 5851 37564
rect 5907 37562 5931 37564
rect 5987 37562 6011 37564
rect 6067 37562 6091 37564
rect 6147 37562 6153 37564
rect 5907 37510 5909 37562
rect 6089 37510 6091 37562
rect 5845 37508 5851 37510
rect 5907 37508 5931 37510
rect 5987 37508 6011 37510
rect 6067 37508 6091 37510
rect 6147 37508 6153 37510
rect 5845 37488 6153 37508
rect 5845 36476 6153 36496
rect 5845 36474 5851 36476
rect 5907 36474 5931 36476
rect 5987 36474 6011 36476
rect 6067 36474 6091 36476
rect 6147 36474 6153 36476
rect 5907 36422 5909 36474
rect 6089 36422 6091 36474
rect 5845 36420 5851 36422
rect 5907 36420 5931 36422
rect 5987 36420 6011 36422
rect 6067 36420 6091 36422
rect 6147 36420 6153 36422
rect 5845 36400 6153 36420
rect 5845 35388 6153 35408
rect 5845 35386 5851 35388
rect 5907 35386 5931 35388
rect 5987 35386 6011 35388
rect 6067 35386 6091 35388
rect 6147 35386 6153 35388
rect 5907 35334 5909 35386
rect 6089 35334 6091 35386
rect 5845 35332 5851 35334
rect 5907 35332 5931 35334
rect 5987 35332 6011 35334
rect 6067 35332 6091 35334
rect 6147 35332 6153 35334
rect 5845 35312 6153 35332
rect 5845 34300 6153 34320
rect 5845 34298 5851 34300
rect 5907 34298 5931 34300
rect 5987 34298 6011 34300
rect 6067 34298 6091 34300
rect 6147 34298 6153 34300
rect 5907 34246 5909 34298
rect 6089 34246 6091 34298
rect 5845 34244 5851 34246
rect 5907 34244 5931 34246
rect 5987 34244 6011 34246
rect 6067 34244 6091 34246
rect 6147 34244 6153 34246
rect 5845 34224 6153 34244
rect 5632 33856 5684 33862
rect 5632 33798 5684 33804
rect 5845 33212 6153 33232
rect 5845 33210 5851 33212
rect 5907 33210 5931 33212
rect 5987 33210 6011 33212
rect 6067 33210 6091 33212
rect 6147 33210 6153 33212
rect 5907 33158 5909 33210
rect 6089 33158 6091 33210
rect 5845 33156 5851 33158
rect 5907 33156 5931 33158
rect 5987 33156 6011 33158
rect 6067 33156 6091 33158
rect 6147 33156 6153 33158
rect 5845 33136 6153 33156
rect 5356 33040 5408 33046
rect 5356 32982 5408 32988
rect 5845 32124 6153 32144
rect 5845 32122 5851 32124
rect 5907 32122 5931 32124
rect 5987 32122 6011 32124
rect 6067 32122 6091 32124
rect 6147 32122 6153 32124
rect 5907 32070 5909 32122
rect 6089 32070 6091 32122
rect 5845 32068 5851 32070
rect 5907 32068 5931 32070
rect 5987 32068 6011 32070
rect 6067 32068 6091 32070
rect 6147 32068 6153 32070
rect 5845 32048 6153 32068
rect 5845 31036 6153 31056
rect 5845 31034 5851 31036
rect 5907 31034 5931 31036
rect 5987 31034 6011 31036
rect 6067 31034 6091 31036
rect 6147 31034 6153 31036
rect 5907 30982 5909 31034
rect 6089 30982 6091 31034
rect 5845 30980 5851 30982
rect 5907 30980 5931 30982
rect 5987 30980 6011 30982
rect 6067 30980 6091 30982
rect 6147 30980 6153 30982
rect 5845 30960 6153 30980
rect 5845 29948 6153 29968
rect 5845 29946 5851 29948
rect 5907 29946 5931 29948
rect 5987 29946 6011 29948
rect 6067 29946 6091 29948
rect 6147 29946 6153 29948
rect 5907 29894 5909 29946
rect 6089 29894 6091 29946
rect 5845 29892 5851 29894
rect 5907 29892 5931 29894
rect 5987 29892 6011 29894
rect 6067 29892 6091 29894
rect 6147 29892 6153 29894
rect 5845 29872 6153 29892
rect 5845 28860 6153 28880
rect 5845 28858 5851 28860
rect 5907 28858 5931 28860
rect 5987 28858 6011 28860
rect 6067 28858 6091 28860
rect 6147 28858 6153 28860
rect 5907 28806 5909 28858
rect 6089 28806 6091 28858
rect 5845 28804 5851 28806
rect 5907 28804 5931 28806
rect 5987 28804 6011 28806
rect 6067 28804 6091 28806
rect 6147 28804 6153 28806
rect 5845 28784 6153 28804
rect 6196 28150 6224 57394
rect 6288 29238 6316 60046
rect 6368 56840 6420 56846
rect 6368 56782 6420 56788
rect 6276 29232 6328 29238
rect 6276 29174 6328 29180
rect 6184 28144 6236 28150
rect 6184 28086 6236 28092
rect 5845 27772 6153 27792
rect 5845 27770 5851 27772
rect 5907 27770 5931 27772
rect 5987 27770 6011 27772
rect 6067 27770 6091 27772
rect 6147 27770 6153 27772
rect 5907 27718 5909 27770
rect 6089 27718 6091 27770
rect 5845 27716 5851 27718
rect 5907 27716 5931 27718
rect 5987 27716 6011 27718
rect 6067 27716 6091 27718
rect 6147 27716 6153 27718
rect 5845 27696 6153 27716
rect 5845 26684 6153 26704
rect 5845 26682 5851 26684
rect 5907 26682 5931 26684
rect 5987 26682 6011 26684
rect 6067 26682 6091 26684
rect 6147 26682 6153 26684
rect 5907 26630 5909 26682
rect 6089 26630 6091 26682
rect 5845 26628 5851 26630
rect 5907 26628 5931 26630
rect 5987 26628 6011 26630
rect 6067 26628 6091 26630
rect 6147 26628 6153 26630
rect 5845 26608 6153 26628
rect 5845 25596 6153 25616
rect 5845 25594 5851 25596
rect 5907 25594 5931 25596
rect 5987 25594 6011 25596
rect 6067 25594 6091 25596
rect 6147 25594 6153 25596
rect 5907 25542 5909 25594
rect 6089 25542 6091 25594
rect 5845 25540 5851 25542
rect 5907 25540 5931 25542
rect 5987 25540 6011 25542
rect 6067 25540 6091 25542
rect 6147 25540 6153 25542
rect 5845 25520 6153 25540
rect 6380 25362 6408 56782
rect 6552 56296 6604 56302
rect 6552 56238 6604 56244
rect 6460 49836 6512 49842
rect 6460 49778 6512 49784
rect 6368 25356 6420 25362
rect 6368 25298 6420 25304
rect 5845 24508 6153 24528
rect 5845 24506 5851 24508
rect 5907 24506 5931 24508
rect 5987 24506 6011 24508
rect 6067 24506 6091 24508
rect 6147 24506 6153 24508
rect 5907 24454 5909 24506
rect 6089 24454 6091 24506
rect 5845 24452 5851 24454
rect 5907 24452 5931 24454
rect 5987 24452 6011 24454
rect 6067 24452 6091 24454
rect 6147 24452 6153 24454
rect 5845 24432 6153 24452
rect 5845 23420 6153 23440
rect 5845 23418 5851 23420
rect 5907 23418 5931 23420
rect 5987 23418 6011 23420
rect 6067 23418 6091 23420
rect 6147 23418 6153 23420
rect 5907 23366 5909 23418
rect 6089 23366 6091 23418
rect 5845 23364 5851 23366
rect 5907 23364 5931 23366
rect 5987 23364 6011 23366
rect 6067 23364 6091 23366
rect 6147 23364 6153 23366
rect 5845 23344 6153 23364
rect 5845 22332 6153 22352
rect 5845 22330 5851 22332
rect 5907 22330 5931 22332
rect 5987 22330 6011 22332
rect 6067 22330 6091 22332
rect 6147 22330 6153 22332
rect 5907 22278 5909 22330
rect 6089 22278 6091 22330
rect 5845 22276 5851 22278
rect 5907 22276 5931 22278
rect 5987 22276 6011 22278
rect 6067 22276 6091 22278
rect 6147 22276 6153 22278
rect 5845 22256 6153 22276
rect 5845 21244 6153 21264
rect 5845 21242 5851 21244
rect 5907 21242 5931 21244
rect 5987 21242 6011 21244
rect 6067 21242 6091 21244
rect 6147 21242 6153 21244
rect 5907 21190 5909 21242
rect 6089 21190 6091 21242
rect 5845 21188 5851 21190
rect 5907 21188 5931 21190
rect 5987 21188 6011 21190
rect 6067 21188 6091 21190
rect 6147 21188 6153 21190
rect 5845 21168 6153 21188
rect 5845 20156 6153 20176
rect 5845 20154 5851 20156
rect 5907 20154 5931 20156
rect 5987 20154 6011 20156
rect 6067 20154 6091 20156
rect 6147 20154 6153 20156
rect 5907 20102 5909 20154
rect 6089 20102 6091 20154
rect 5845 20100 5851 20102
rect 5907 20100 5931 20102
rect 5987 20100 6011 20102
rect 6067 20100 6091 20102
rect 6147 20100 6153 20102
rect 5845 20080 6153 20100
rect 5845 19068 6153 19088
rect 5845 19066 5851 19068
rect 5907 19066 5931 19068
rect 5987 19066 6011 19068
rect 6067 19066 6091 19068
rect 6147 19066 6153 19068
rect 5907 19014 5909 19066
rect 6089 19014 6091 19066
rect 5845 19012 5851 19014
rect 5907 19012 5931 19014
rect 5987 19012 6011 19014
rect 6067 19012 6091 19014
rect 6147 19012 6153 19014
rect 5845 18992 6153 19012
rect 5845 17980 6153 18000
rect 5845 17978 5851 17980
rect 5907 17978 5931 17980
rect 5987 17978 6011 17980
rect 6067 17978 6091 17980
rect 6147 17978 6153 17980
rect 5907 17926 5909 17978
rect 6089 17926 6091 17978
rect 5845 17924 5851 17926
rect 5907 17924 5931 17926
rect 5987 17924 6011 17926
rect 6067 17924 6091 17926
rect 6147 17924 6153 17926
rect 5845 17904 6153 17924
rect 6472 17882 6500 49778
rect 6564 23594 6592 56238
rect 6644 51876 6696 51882
rect 6644 51818 6696 51824
rect 6552 23588 6604 23594
rect 6552 23530 6604 23536
rect 6656 23050 6684 51818
rect 6748 51074 6776 63718
rect 6748 51046 6868 51074
rect 6736 50788 6788 50794
rect 6736 50730 6788 50736
rect 6748 46442 6776 50730
rect 6840 48793 6868 51046
rect 6826 48784 6882 48793
rect 6826 48719 6882 48728
rect 6828 48680 6880 48686
rect 6828 48622 6880 48628
rect 6736 46436 6788 46442
rect 6736 46378 6788 46384
rect 6734 46336 6790 46345
rect 6734 46271 6790 46280
rect 6748 41614 6776 46271
rect 6736 41608 6788 41614
rect 6736 41550 6788 41556
rect 6644 23044 6696 23050
rect 6644 22986 6696 22992
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 5845 16892 6153 16912
rect 5845 16890 5851 16892
rect 5907 16890 5931 16892
rect 5987 16890 6011 16892
rect 6067 16890 6091 16892
rect 6147 16890 6153 16892
rect 5907 16838 5909 16890
rect 6089 16838 6091 16890
rect 5845 16836 5851 16838
rect 5907 16836 5931 16838
rect 5987 16836 6011 16838
rect 6067 16836 6091 16838
rect 6147 16836 6153 16838
rect 5845 16816 6153 16836
rect 5845 15804 6153 15824
rect 5845 15802 5851 15804
rect 5907 15802 5931 15804
rect 5987 15802 6011 15804
rect 6067 15802 6091 15804
rect 6147 15802 6153 15804
rect 5907 15750 5909 15802
rect 6089 15750 6091 15802
rect 5845 15748 5851 15750
rect 5907 15748 5931 15750
rect 5987 15748 6011 15750
rect 6067 15748 6091 15750
rect 6147 15748 6153 15750
rect 5845 15728 6153 15748
rect 5845 14716 6153 14736
rect 5845 14714 5851 14716
rect 5907 14714 5931 14716
rect 5987 14714 6011 14716
rect 6067 14714 6091 14716
rect 6147 14714 6153 14716
rect 5907 14662 5909 14714
rect 6089 14662 6091 14714
rect 5845 14660 5851 14662
rect 5907 14660 5931 14662
rect 5987 14660 6011 14662
rect 6067 14660 6091 14662
rect 6147 14660 6153 14662
rect 5845 14640 6153 14660
rect 5845 13628 6153 13648
rect 5845 13626 5851 13628
rect 5907 13626 5931 13628
rect 5987 13626 6011 13628
rect 6067 13626 6091 13628
rect 6147 13626 6153 13628
rect 5907 13574 5909 13626
rect 6089 13574 6091 13626
rect 5845 13572 5851 13574
rect 5907 13572 5931 13574
rect 5987 13572 6011 13574
rect 6067 13572 6091 13574
rect 6147 13572 6153 13574
rect 5845 13552 6153 13572
rect 5845 12540 6153 12560
rect 5845 12538 5851 12540
rect 5907 12538 5931 12540
rect 5987 12538 6011 12540
rect 6067 12538 6091 12540
rect 6147 12538 6153 12540
rect 5907 12486 5909 12538
rect 6089 12486 6091 12538
rect 5845 12484 5851 12486
rect 5907 12484 5931 12486
rect 5987 12484 6011 12486
rect 6067 12484 6091 12486
rect 6147 12484 6153 12486
rect 5845 12464 6153 12484
rect 5845 11452 6153 11472
rect 5845 11450 5851 11452
rect 5907 11450 5931 11452
rect 5987 11450 6011 11452
rect 6067 11450 6091 11452
rect 6147 11450 6153 11452
rect 5907 11398 5909 11450
rect 6089 11398 6091 11450
rect 5845 11396 5851 11398
rect 5907 11396 5931 11398
rect 5987 11396 6011 11398
rect 6067 11396 6091 11398
rect 6147 11396 6153 11398
rect 5845 11376 6153 11396
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4632 10062 4660 10542
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4213 9820 4521 9840
rect 4213 9818 4219 9820
rect 4275 9818 4299 9820
rect 4355 9818 4379 9820
rect 4435 9818 4459 9820
rect 4515 9818 4521 9820
rect 4275 9766 4277 9818
rect 4457 9766 4459 9818
rect 4213 9764 4219 9766
rect 4275 9764 4299 9766
rect 4355 9764 4379 9766
rect 4435 9764 4459 9766
rect 4515 9764 4521 9766
rect 4213 9744 4521 9764
rect 4632 9586 4660 9998
rect 4908 9586 4936 10610
rect 5845 10364 6153 10384
rect 5845 10362 5851 10364
rect 5907 10362 5931 10364
rect 5987 10362 6011 10364
rect 6067 10362 6091 10364
rect 6147 10362 6153 10364
rect 5907 10310 5909 10362
rect 6089 10310 6091 10362
rect 5845 10308 5851 10310
rect 5907 10308 5931 10310
rect 5987 10308 6011 10310
rect 6067 10308 6091 10310
rect 6147 10308 6153 10310
rect 5845 10288 6153 10308
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4213 8732 4521 8752
rect 4213 8730 4219 8732
rect 4275 8730 4299 8732
rect 4355 8730 4379 8732
rect 4435 8730 4459 8732
rect 4515 8730 4521 8732
rect 4275 8678 4277 8730
rect 4457 8678 4459 8730
rect 4213 8676 4219 8678
rect 4275 8676 4299 8678
rect 4355 8676 4379 8678
rect 4435 8676 4459 8678
rect 4515 8676 4521 8678
rect 4213 8656 4521 8676
rect 4632 7886 4660 9522
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1216 4140 1268 4146
rect 1216 4082 1268 4088
rect 1228 3369 1256 4082
rect 1412 3777 1440 4558
rect 1398 3768 1454 3777
rect 1398 3703 1454 3712
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1214 3360 1270 3369
rect 1214 3295 1270 3304
rect 1320 2825 1348 3470
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1306 2816 1362 2825
rect 1306 2751 1362 2760
rect 1308 2440 1360 2446
rect 1412 2417 1440 2994
rect 1504 2650 1532 5646
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 3194 1624 5170
rect 1688 3738 1716 6258
rect 2582 6012 2890 6032
rect 2582 6010 2588 6012
rect 2644 6010 2668 6012
rect 2724 6010 2748 6012
rect 2804 6010 2828 6012
rect 2884 6010 2890 6012
rect 2644 5958 2646 6010
rect 2826 5958 2828 6010
rect 2582 5956 2588 5958
rect 2644 5956 2668 5958
rect 2724 5956 2748 5958
rect 2804 5956 2828 5958
rect 2884 5956 2890 5958
rect 2582 5936 2890 5956
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 2148 2650 2176 5646
rect 2976 5370 3004 6734
rect 3896 6458 3924 7822
rect 4213 7644 4521 7664
rect 4213 7642 4219 7644
rect 4275 7642 4299 7644
rect 4355 7642 4379 7644
rect 4435 7642 4459 7644
rect 4515 7642 4521 7644
rect 4275 7590 4277 7642
rect 4457 7590 4459 7642
rect 4213 7588 4219 7590
rect 4275 7588 4299 7590
rect 4355 7588 4379 7590
rect 4435 7588 4459 7590
rect 4515 7588 4521 7590
rect 4213 7568 4521 7588
rect 5092 6798 5120 9454
rect 5845 9276 6153 9296
rect 5845 9274 5851 9276
rect 5907 9274 5931 9276
rect 5987 9274 6011 9276
rect 6067 9274 6091 9276
rect 6147 9274 6153 9276
rect 5907 9222 5909 9274
rect 6089 9222 6091 9274
rect 5845 9220 5851 9222
rect 5907 9220 5931 9222
rect 5987 9220 6011 9222
rect 6067 9220 6091 9222
rect 6147 9220 6153 9222
rect 5845 9200 6153 9220
rect 5845 8188 6153 8208
rect 5845 8186 5851 8188
rect 5907 8186 5931 8188
rect 5987 8186 6011 8188
rect 6067 8186 6091 8188
rect 6147 8186 6153 8188
rect 5907 8134 5909 8186
rect 6089 8134 6091 8186
rect 5845 8132 5851 8134
rect 5907 8132 5931 8134
rect 5987 8132 6011 8134
rect 6067 8132 6091 8134
rect 6147 8132 6153 8134
rect 5845 8112 6153 8132
rect 5845 7100 6153 7120
rect 5845 7098 5851 7100
rect 5907 7098 5931 7100
rect 5987 7098 6011 7100
rect 6067 7098 6091 7100
rect 6147 7098 6153 7100
rect 5907 7046 5909 7098
rect 6089 7046 6091 7098
rect 5845 7044 5851 7046
rect 5907 7044 5931 7046
rect 5987 7044 6011 7046
rect 6067 7044 6091 7046
rect 6147 7044 6153 7046
rect 5845 7024 6153 7044
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 4213 6556 4521 6576
rect 4213 6554 4219 6556
rect 4275 6554 4299 6556
rect 4355 6554 4379 6556
rect 4435 6554 4459 6556
rect 4515 6554 4521 6556
rect 4275 6502 4277 6554
rect 4457 6502 4459 6554
rect 4213 6500 4219 6502
rect 4275 6500 4299 6502
rect 4355 6500 4379 6502
rect 4435 6500 4459 6502
rect 4515 6500 4521 6502
rect 4213 6480 4521 6500
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 5092 6322 5120 6734
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2582 4924 2890 4944
rect 2582 4922 2588 4924
rect 2644 4922 2668 4924
rect 2724 4922 2748 4924
rect 2804 4922 2828 4924
rect 2884 4922 2890 4924
rect 2644 4870 2646 4922
rect 2826 4870 2828 4922
rect 2582 4868 2588 4870
rect 2644 4868 2668 4870
rect 2724 4868 2748 4870
rect 2804 4868 2828 4870
rect 2884 4868 2890 4870
rect 2582 4848 2890 4868
rect 2976 4010 3004 5170
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2582 3836 2890 3856
rect 2582 3834 2588 3836
rect 2644 3834 2668 3836
rect 2724 3834 2748 3836
rect 2804 3834 2828 3836
rect 2884 3834 2890 3836
rect 2644 3782 2646 3834
rect 2826 3782 2828 3834
rect 2582 3780 2588 3782
rect 2644 3780 2668 3782
rect 2724 3780 2748 3782
rect 2804 3780 2828 3782
rect 2884 3780 2890 3782
rect 2582 3760 2890 3780
rect 3068 2774 3096 5646
rect 3160 4826 3188 6258
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3896 5914 3924 6122
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 5092 5710 5120 6258
rect 6840 6186 6868 48622
rect 6932 42362 6960 67798
rect 7477 67484 7785 67504
rect 7477 67482 7483 67484
rect 7539 67482 7563 67484
rect 7619 67482 7643 67484
rect 7699 67482 7723 67484
rect 7779 67482 7785 67484
rect 7539 67430 7541 67482
rect 7721 67430 7723 67482
rect 7477 67428 7483 67430
rect 7539 67428 7563 67430
rect 7619 67428 7643 67430
rect 7699 67428 7723 67430
rect 7779 67428 7785 67430
rect 7477 67408 7785 67428
rect 7477 66396 7785 66416
rect 7477 66394 7483 66396
rect 7539 66394 7563 66396
rect 7619 66394 7643 66396
rect 7699 66394 7723 66396
rect 7779 66394 7785 66396
rect 7539 66342 7541 66394
rect 7721 66342 7723 66394
rect 7477 66340 7483 66342
rect 7539 66340 7563 66342
rect 7619 66340 7643 66342
rect 7699 66340 7723 66342
rect 7779 66340 7785 66342
rect 7477 66320 7785 66340
rect 7477 65308 7785 65328
rect 7477 65306 7483 65308
rect 7539 65306 7563 65308
rect 7619 65306 7643 65308
rect 7699 65306 7723 65308
rect 7779 65306 7785 65308
rect 7539 65254 7541 65306
rect 7721 65254 7723 65306
rect 7477 65252 7483 65254
rect 7539 65252 7563 65254
rect 7619 65252 7643 65254
rect 7699 65252 7723 65254
rect 7779 65252 7785 65254
rect 7477 65232 7785 65252
rect 7477 64220 7785 64240
rect 7477 64218 7483 64220
rect 7539 64218 7563 64220
rect 7619 64218 7643 64220
rect 7699 64218 7723 64220
rect 7779 64218 7785 64220
rect 7539 64166 7541 64218
rect 7721 64166 7723 64218
rect 7477 64164 7483 64166
rect 7539 64164 7563 64166
rect 7619 64164 7643 64166
rect 7699 64164 7723 64166
rect 7779 64164 7785 64166
rect 7477 64144 7785 64164
rect 7380 63300 7432 63306
rect 7380 63242 7432 63248
rect 7288 62144 7340 62150
rect 7288 62086 7340 62092
rect 7012 54188 7064 54194
rect 7012 54130 7064 54136
rect 6920 42356 6972 42362
rect 6920 42298 6972 42304
rect 7024 19990 7052 54130
rect 7104 54120 7156 54126
rect 7104 54062 7156 54068
rect 7116 20058 7144 54062
rect 7196 53508 7248 53514
rect 7196 53450 7248 53456
rect 7208 20398 7236 53450
rect 7300 33930 7328 62086
rect 7392 38486 7420 63242
rect 7477 63132 7785 63152
rect 7477 63130 7483 63132
rect 7539 63130 7563 63132
rect 7619 63130 7643 63132
rect 7699 63130 7723 63132
rect 7779 63130 7785 63132
rect 7539 63078 7541 63130
rect 7721 63078 7723 63130
rect 7477 63076 7483 63078
rect 7539 63076 7563 63078
rect 7619 63076 7643 63078
rect 7699 63076 7723 63078
rect 7779 63076 7785 63078
rect 7477 63056 7785 63076
rect 7477 62044 7785 62064
rect 7477 62042 7483 62044
rect 7539 62042 7563 62044
rect 7619 62042 7643 62044
rect 7699 62042 7723 62044
rect 7779 62042 7785 62044
rect 7539 61990 7541 62042
rect 7721 61990 7723 62042
rect 7477 61988 7483 61990
rect 7539 61988 7563 61990
rect 7619 61988 7643 61990
rect 7699 61988 7723 61990
rect 7779 61988 7785 61990
rect 7477 61968 7785 61988
rect 7477 60956 7785 60976
rect 7477 60954 7483 60956
rect 7539 60954 7563 60956
rect 7619 60954 7643 60956
rect 7699 60954 7723 60956
rect 7779 60954 7785 60956
rect 7539 60902 7541 60954
rect 7721 60902 7723 60954
rect 7477 60900 7483 60902
rect 7539 60900 7563 60902
rect 7619 60900 7643 60902
rect 7699 60900 7723 60902
rect 7779 60900 7785 60902
rect 7477 60880 7785 60900
rect 7477 59868 7785 59888
rect 7477 59866 7483 59868
rect 7539 59866 7563 59868
rect 7619 59866 7643 59868
rect 7699 59866 7723 59868
rect 7779 59866 7785 59868
rect 7539 59814 7541 59866
rect 7721 59814 7723 59866
rect 7477 59812 7483 59814
rect 7539 59812 7563 59814
rect 7619 59812 7643 59814
rect 7699 59812 7723 59814
rect 7779 59812 7785 59814
rect 7477 59792 7785 59812
rect 7477 58780 7785 58800
rect 7477 58778 7483 58780
rect 7539 58778 7563 58780
rect 7619 58778 7643 58780
rect 7699 58778 7723 58780
rect 7779 58778 7785 58780
rect 7539 58726 7541 58778
rect 7721 58726 7723 58778
rect 7477 58724 7483 58726
rect 7539 58724 7563 58726
rect 7619 58724 7643 58726
rect 7699 58724 7723 58726
rect 7779 58724 7785 58726
rect 7477 58704 7785 58724
rect 7477 57692 7785 57712
rect 7477 57690 7483 57692
rect 7539 57690 7563 57692
rect 7619 57690 7643 57692
rect 7699 57690 7723 57692
rect 7779 57690 7785 57692
rect 7539 57638 7541 57690
rect 7721 57638 7723 57690
rect 7477 57636 7483 57638
rect 7539 57636 7563 57638
rect 7619 57636 7643 57638
rect 7699 57636 7723 57638
rect 7779 57636 7785 57638
rect 7477 57616 7785 57636
rect 7477 56604 7785 56624
rect 7477 56602 7483 56604
rect 7539 56602 7563 56604
rect 7619 56602 7643 56604
rect 7699 56602 7723 56604
rect 7779 56602 7785 56604
rect 7539 56550 7541 56602
rect 7721 56550 7723 56602
rect 7477 56548 7483 56550
rect 7539 56548 7563 56550
rect 7619 56548 7643 56550
rect 7699 56548 7723 56550
rect 7779 56548 7785 56550
rect 7477 56528 7785 56548
rect 7477 55516 7785 55536
rect 7477 55514 7483 55516
rect 7539 55514 7563 55516
rect 7619 55514 7643 55516
rect 7699 55514 7723 55516
rect 7779 55514 7785 55516
rect 7539 55462 7541 55514
rect 7721 55462 7723 55514
rect 7477 55460 7483 55462
rect 7539 55460 7563 55462
rect 7619 55460 7643 55462
rect 7699 55460 7723 55462
rect 7779 55460 7785 55462
rect 7477 55440 7785 55460
rect 7840 55344 7892 55350
rect 7840 55286 7892 55292
rect 7477 54428 7785 54448
rect 7477 54426 7483 54428
rect 7539 54426 7563 54428
rect 7619 54426 7643 54428
rect 7699 54426 7723 54428
rect 7779 54426 7785 54428
rect 7539 54374 7541 54426
rect 7721 54374 7723 54426
rect 7477 54372 7483 54374
rect 7539 54372 7563 54374
rect 7619 54372 7643 54374
rect 7699 54372 7723 54374
rect 7779 54372 7785 54374
rect 7477 54352 7785 54372
rect 7477 53340 7785 53360
rect 7477 53338 7483 53340
rect 7539 53338 7563 53340
rect 7619 53338 7643 53340
rect 7699 53338 7723 53340
rect 7779 53338 7785 53340
rect 7539 53286 7541 53338
rect 7721 53286 7723 53338
rect 7477 53284 7483 53286
rect 7539 53284 7563 53286
rect 7619 53284 7643 53286
rect 7699 53284 7723 53286
rect 7779 53284 7785 53286
rect 7477 53264 7785 53284
rect 7477 52252 7785 52272
rect 7477 52250 7483 52252
rect 7539 52250 7563 52252
rect 7619 52250 7643 52252
rect 7699 52250 7723 52252
rect 7779 52250 7785 52252
rect 7539 52198 7541 52250
rect 7721 52198 7723 52250
rect 7477 52196 7483 52198
rect 7539 52196 7563 52198
rect 7619 52196 7643 52198
rect 7699 52196 7723 52198
rect 7779 52196 7785 52198
rect 7477 52176 7785 52196
rect 7477 51164 7785 51184
rect 7477 51162 7483 51164
rect 7539 51162 7563 51164
rect 7619 51162 7643 51164
rect 7699 51162 7723 51164
rect 7779 51162 7785 51164
rect 7539 51110 7541 51162
rect 7721 51110 7723 51162
rect 7477 51108 7483 51110
rect 7539 51108 7563 51110
rect 7619 51108 7643 51110
rect 7699 51108 7723 51110
rect 7779 51108 7785 51110
rect 7477 51088 7785 51108
rect 7477 50076 7785 50096
rect 7477 50074 7483 50076
rect 7539 50074 7563 50076
rect 7619 50074 7643 50076
rect 7699 50074 7723 50076
rect 7779 50074 7785 50076
rect 7539 50022 7541 50074
rect 7721 50022 7723 50074
rect 7477 50020 7483 50022
rect 7539 50020 7563 50022
rect 7619 50020 7643 50022
rect 7699 50020 7723 50022
rect 7779 50020 7785 50022
rect 7477 50000 7785 50020
rect 7477 48988 7785 49008
rect 7477 48986 7483 48988
rect 7539 48986 7563 48988
rect 7619 48986 7643 48988
rect 7699 48986 7723 48988
rect 7779 48986 7785 48988
rect 7539 48934 7541 48986
rect 7721 48934 7723 48986
rect 7477 48932 7483 48934
rect 7539 48932 7563 48934
rect 7619 48932 7643 48934
rect 7699 48932 7723 48934
rect 7779 48932 7785 48934
rect 7477 48912 7785 48932
rect 7477 47900 7785 47920
rect 7477 47898 7483 47900
rect 7539 47898 7563 47900
rect 7619 47898 7643 47900
rect 7699 47898 7723 47900
rect 7779 47898 7785 47900
rect 7539 47846 7541 47898
rect 7721 47846 7723 47898
rect 7477 47844 7483 47846
rect 7539 47844 7563 47846
rect 7619 47844 7643 47846
rect 7699 47844 7723 47846
rect 7779 47844 7785 47846
rect 7477 47824 7785 47844
rect 7477 46812 7785 46832
rect 7477 46810 7483 46812
rect 7539 46810 7563 46812
rect 7619 46810 7643 46812
rect 7699 46810 7723 46812
rect 7779 46810 7785 46812
rect 7539 46758 7541 46810
rect 7721 46758 7723 46810
rect 7477 46756 7483 46758
rect 7539 46756 7563 46758
rect 7619 46756 7643 46758
rect 7699 46756 7723 46758
rect 7779 46756 7785 46758
rect 7477 46736 7785 46756
rect 7477 45724 7785 45744
rect 7477 45722 7483 45724
rect 7539 45722 7563 45724
rect 7619 45722 7643 45724
rect 7699 45722 7723 45724
rect 7779 45722 7785 45724
rect 7539 45670 7541 45722
rect 7721 45670 7723 45722
rect 7477 45668 7483 45670
rect 7539 45668 7563 45670
rect 7619 45668 7643 45670
rect 7699 45668 7723 45670
rect 7779 45668 7785 45670
rect 7477 45648 7785 45668
rect 7477 44636 7785 44656
rect 7477 44634 7483 44636
rect 7539 44634 7563 44636
rect 7619 44634 7643 44636
rect 7699 44634 7723 44636
rect 7779 44634 7785 44636
rect 7539 44582 7541 44634
rect 7721 44582 7723 44634
rect 7477 44580 7483 44582
rect 7539 44580 7563 44582
rect 7619 44580 7643 44582
rect 7699 44580 7723 44582
rect 7779 44580 7785 44582
rect 7477 44560 7785 44580
rect 7477 43548 7785 43568
rect 7477 43546 7483 43548
rect 7539 43546 7563 43548
rect 7619 43546 7643 43548
rect 7699 43546 7723 43548
rect 7779 43546 7785 43548
rect 7539 43494 7541 43546
rect 7721 43494 7723 43546
rect 7477 43492 7483 43494
rect 7539 43492 7563 43494
rect 7619 43492 7643 43494
rect 7699 43492 7723 43494
rect 7779 43492 7785 43494
rect 7477 43472 7785 43492
rect 7477 42460 7785 42480
rect 7477 42458 7483 42460
rect 7539 42458 7563 42460
rect 7619 42458 7643 42460
rect 7699 42458 7723 42460
rect 7779 42458 7785 42460
rect 7539 42406 7541 42458
rect 7721 42406 7723 42458
rect 7477 42404 7483 42406
rect 7539 42404 7563 42406
rect 7619 42404 7643 42406
rect 7699 42404 7723 42406
rect 7779 42404 7785 42406
rect 7477 42384 7785 42404
rect 7477 41372 7785 41392
rect 7477 41370 7483 41372
rect 7539 41370 7563 41372
rect 7619 41370 7643 41372
rect 7699 41370 7723 41372
rect 7779 41370 7785 41372
rect 7539 41318 7541 41370
rect 7721 41318 7723 41370
rect 7477 41316 7483 41318
rect 7539 41316 7563 41318
rect 7619 41316 7643 41318
rect 7699 41316 7723 41318
rect 7779 41316 7785 41318
rect 7477 41296 7785 41316
rect 7477 40284 7785 40304
rect 7477 40282 7483 40284
rect 7539 40282 7563 40284
rect 7619 40282 7643 40284
rect 7699 40282 7723 40284
rect 7779 40282 7785 40284
rect 7539 40230 7541 40282
rect 7721 40230 7723 40282
rect 7477 40228 7483 40230
rect 7539 40228 7563 40230
rect 7619 40228 7643 40230
rect 7699 40228 7723 40230
rect 7779 40228 7785 40230
rect 7477 40208 7785 40228
rect 7477 39196 7785 39216
rect 7477 39194 7483 39196
rect 7539 39194 7563 39196
rect 7619 39194 7643 39196
rect 7699 39194 7723 39196
rect 7779 39194 7785 39196
rect 7539 39142 7541 39194
rect 7721 39142 7723 39194
rect 7477 39140 7483 39142
rect 7539 39140 7563 39142
rect 7619 39140 7643 39142
rect 7699 39140 7723 39142
rect 7779 39140 7785 39142
rect 7477 39120 7785 39140
rect 7380 38480 7432 38486
rect 7380 38422 7432 38428
rect 7477 38108 7785 38128
rect 7477 38106 7483 38108
rect 7539 38106 7563 38108
rect 7619 38106 7643 38108
rect 7699 38106 7723 38108
rect 7779 38106 7785 38108
rect 7539 38054 7541 38106
rect 7721 38054 7723 38106
rect 7477 38052 7483 38054
rect 7539 38052 7563 38054
rect 7619 38052 7643 38054
rect 7699 38052 7723 38054
rect 7779 38052 7785 38054
rect 7477 38032 7785 38052
rect 7477 37020 7785 37040
rect 7477 37018 7483 37020
rect 7539 37018 7563 37020
rect 7619 37018 7643 37020
rect 7699 37018 7723 37020
rect 7779 37018 7785 37020
rect 7539 36966 7541 37018
rect 7721 36966 7723 37018
rect 7477 36964 7483 36966
rect 7539 36964 7563 36966
rect 7619 36964 7643 36966
rect 7699 36964 7723 36966
rect 7779 36964 7785 36966
rect 7477 36944 7785 36964
rect 7477 35932 7785 35952
rect 7477 35930 7483 35932
rect 7539 35930 7563 35932
rect 7619 35930 7643 35932
rect 7699 35930 7723 35932
rect 7779 35930 7785 35932
rect 7539 35878 7541 35930
rect 7721 35878 7723 35930
rect 7477 35876 7483 35878
rect 7539 35876 7563 35878
rect 7619 35876 7643 35878
rect 7699 35876 7723 35878
rect 7779 35876 7785 35878
rect 7477 35856 7785 35876
rect 7477 34844 7785 34864
rect 7477 34842 7483 34844
rect 7539 34842 7563 34844
rect 7619 34842 7643 34844
rect 7699 34842 7723 34844
rect 7779 34842 7785 34844
rect 7539 34790 7541 34842
rect 7721 34790 7723 34842
rect 7477 34788 7483 34790
rect 7539 34788 7563 34790
rect 7619 34788 7643 34790
rect 7699 34788 7723 34790
rect 7779 34788 7785 34790
rect 7477 34768 7785 34788
rect 7288 33924 7340 33930
rect 7288 33866 7340 33872
rect 7477 33756 7785 33776
rect 7477 33754 7483 33756
rect 7539 33754 7563 33756
rect 7619 33754 7643 33756
rect 7699 33754 7723 33756
rect 7779 33754 7785 33756
rect 7539 33702 7541 33754
rect 7721 33702 7723 33754
rect 7477 33700 7483 33702
rect 7539 33700 7563 33702
rect 7619 33700 7643 33702
rect 7699 33700 7723 33702
rect 7779 33700 7785 33702
rect 7477 33680 7785 33700
rect 7477 32668 7785 32688
rect 7477 32666 7483 32668
rect 7539 32666 7563 32668
rect 7619 32666 7643 32668
rect 7699 32666 7723 32668
rect 7779 32666 7785 32668
rect 7539 32614 7541 32666
rect 7721 32614 7723 32666
rect 7477 32612 7483 32614
rect 7539 32612 7563 32614
rect 7619 32612 7643 32614
rect 7699 32612 7723 32614
rect 7779 32612 7785 32614
rect 7477 32592 7785 32612
rect 7477 31580 7785 31600
rect 7477 31578 7483 31580
rect 7539 31578 7563 31580
rect 7619 31578 7643 31580
rect 7699 31578 7723 31580
rect 7779 31578 7785 31580
rect 7539 31526 7541 31578
rect 7721 31526 7723 31578
rect 7477 31524 7483 31526
rect 7539 31524 7563 31526
rect 7619 31524 7643 31526
rect 7699 31524 7723 31526
rect 7779 31524 7785 31526
rect 7477 31504 7785 31524
rect 7477 30492 7785 30512
rect 7477 30490 7483 30492
rect 7539 30490 7563 30492
rect 7619 30490 7643 30492
rect 7699 30490 7723 30492
rect 7779 30490 7785 30492
rect 7539 30438 7541 30490
rect 7721 30438 7723 30490
rect 7477 30436 7483 30438
rect 7539 30436 7563 30438
rect 7619 30436 7643 30438
rect 7699 30436 7723 30438
rect 7779 30436 7785 30438
rect 7477 30416 7785 30436
rect 7477 29404 7785 29424
rect 7477 29402 7483 29404
rect 7539 29402 7563 29404
rect 7619 29402 7643 29404
rect 7699 29402 7723 29404
rect 7779 29402 7785 29404
rect 7539 29350 7541 29402
rect 7721 29350 7723 29402
rect 7477 29348 7483 29350
rect 7539 29348 7563 29350
rect 7619 29348 7643 29350
rect 7699 29348 7723 29350
rect 7779 29348 7785 29350
rect 7477 29328 7785 29348
rect 7477 28316 7785 28336
rect 7477 28314 7483 28316
rect 7539 28314 7563 28316
rect 7619 28314 7643 28316
rect 7699 28314 7723 28316
rect 7779 28314 7785 28316
rect 7539 28262 7541 28314
rect 7721 28262 7723 28314
rect 7477 28260 7483 28262
rect 7539 28260 7563 28262
rect 7619 28260 7643 28262
rect 7699 28260 7723 28262
rect 7779 28260 7785 28262
rect 7477 28240 7785 28260
rect 7477 27228 7785 27248
rect 7477 27226 7483 27228
rect 7539 27226 7563 27228
rect 7619 27226 7643 27228
rect 7699 27226 7723 27228
rect 7779 27226 7785 27228
rect 7539 27174 7541 27226
rect 7721 27174 7723 27226
rect 7477 27172 7483 27174
rect 7539 27172 7563 27174
rect 7619 27172 7643 27174
rect 7699 27172 7723 27174
rect 7779 27172 7785 27174
rect 7477 27152 7785 27172
rect 7477 26140 7785 26160
rect 7477 26138 7483 26140
rect 7539 26138 7563 26140
rect 7619 26138 7643 26140
rect 7699 26138 7723 26140
rect 7779 26138 7785 26140
rect 7539 26086 7541 26138
rect 7721 26086 7723 26138
rect 7477 26084 7483 26086
rect 7539 26084 7563 26086
rect 7619 26084 7643 26086
rect 7699 26084 7723 26086
rect 7779 26084 7785 26086
rect 7477 26064 7785 26084
rect 7477 25052 7785 25072
rect 7477 25050 7483 25052
rect 7539 25050 7563 25052
rect 7619 25050 7643 25052
rect 7699 25050 7723 25052
rect 7779 25050 7785 25052
rect 7539 24998 7541 25050
rect 7721 24998 7723 25050
rect 7477 24996 7483 24998
rect 7539 24996 7563 24998
rect 7619 24996 7643 24998
rect 7699 24996 7723 24998
rect 7779 24996 7785 24998
rect 7477 24976 7785 24996
rect 7477 23964 7785 23984
rect 7477 23962 7483 23964
rect 7539 23962 7563 23964
rect 7619 23962 7643 23964
rect 7699 23962 7723 23964
rect 7779 23962 7785 23964
rect 7539 23910 7541 23962
rect 7721 23910 7723 23962
rect 7477 23908 7483 23910
rect 7539 23908 7563 23910
rect 7619 23908 7643 23910
rect 7699 23908 7723 23910
rect 7779 23908 7785 23910
rect 7477 23888 7785 23908
rect 7477 22876 7785 22896
rect 7477 22874 7483 22876
rect 7539 22874 7563 22876
rect 7619 22874 7643 22876
rect 7699 22874 7723 22876
rect 7779 22874 7785 22876
rect 7539 22822 7541 22874
rect 7721 22822 7723 22874
rect 7477 22820 7483 22822
rect 7539 22820 7563 22822
rect 7619 22820 7643 22822
rect 7699 22820 7723 22822
rect 7779 22820 7785 22822
rect 7477 22800 7785 22820
rect 7477 21788 7785 21808
rect 7477 21786 7483 21788
rect 7539 21786 7563 21788
rect 7619 21786 7643 21788
rect 7699 21786 7723 21788
rect 7779 21786 7785 21788
rect 7539 21734 7541 21786
rect 7721 21734 7723 21786
rect 7477 21732 7483 21734
rect 7539 21732 7563 21734
rect 7619 21732 7643 21734
rect 7699 21732 7723 21734
rect 7779 21732 7785 21734
rect 7477 21712 7785 21732
rect 7477 20700 7785 20720
rect 7477 20698 7483 20700
rect 7539 20698 7563 20700
rect 7619 20698 7643 20700
rect 7699 20698 7723 20700
rect 7779 20698 7785 20700
rect 7539 20646 7541 20698
rect 7721 20646 7723 20698
rect 7477 20644 7483 20646
rect 7539 20644 7563 20646
rect 7619 20644 7643 20646
rect 7699 20644 7723 20646
rect 7779 20644 7785 20646
rect 7477 20624 7785 20644
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7012 19984 7064 19990
rect 7012 19926 7064 19932
rect 7477 19612 7785 19632
rect 7477 19610 7483 19612
rect 7539 19610 7563 19612
rect 7619 19610 7643 19612
rect 7699 19610 7723 19612
rect 7779 19610 7785 19612
rect 7539 19558 7541 19610
rect 7721 19558 7723 19610
rect 7477 19556 7483 19558
rect 7539 19556 7563 19558
rect 7619 19556 7643 19558
rect 7699 19556 7723 19558
rect 7779 19556 7785 19558
rect 7477 19536 7785 19556
rect 7852 18698 7880 55286
rect 8312 46918 8340 74326
rect 9784 74186 9812 76230
rect 9968 75342 9996 76774
rect 10140 76424 10192 76430
rect 10140 76366 10192 76372
rect 10152 76129 10180 76366
rect 10138 76120 10194 76129
rect 10138 76055 10194 76064
rect 9956 75336 10008 75342
rect 9956 75278 10008 75284
rect 10140 75336 10192 75342
rect 10140 75278 10192 75284
rect 9864 75200 9916 75206
rect 9864 75142 9916 75148
rect 9772 74180 9824 74186
rect 9772 74122 9824 74128
rect 9876 73846 9904 75142
rect 10152 75041 10180 75278
rect 10138 75032 10194 75041
rect 10138 74967 10194 74976
rect 10140 74248 10192 74254
rect 10140 74190 10192 74196
rect 9956 74112 10008 74118
rect 9956 74054 10008 74060
rect 9864 73840 9916 73846
rect 9864 73782 9916 73788
rect 9109 73468 9417 73488
rect 9109 73466 9115 73468
rect 9171 73466 9195 73468
rect 9251 73466 9275 73468
rect 9331 73466 9355 73468
rect 9411 73466 9417 73468
rect 9171 73414 9173 73466
rect 9353 73414 9355 73466
rect 9109 73412 9115 73414
rect 9171 73412 9195 73414
rect 9251 73412 9275 73414
rect 9331 73412 9355 73414
rect 9411 73412 9417 73414
rect 9109 73392 9417 73412
rect 9968 73166 9996 74054
rect 10152 73953 10180 74190
rect 10138 73944 10194 73953
rect 10138 73879 10194 73888
rect 9956 73160 10008 73166
rect 9956 73102 10008 73108
rect 10140 73160 10192 73166
rect 10140 73102 10192 73108
rect 8392 73024 8444 73030
rect 8392 72966 8444 72972
rect 8404 72010 8432 72966
rect 10152 72729 10180 73102
rect 10138 72720 10194 72729
rect 10138 72655 10194 72664
rect 9109 72380 9417 72400
rect 9109 72378 9115 72380
rect 9171 72378 9195 72380
rect 9251 72378 9275 72380
rect 9331 72378 9355 72380
rect 9411 72378 9417 72380
rect 9171 72326 9173 72378
rect 9353 72326 9355 72378
rect 9109 72324 9115 72326
rect 9171 72324 9195 72326
rect 9251 72324 9275 72326
rect 9331 72324 9355 72326
rect 9411 72324 9417 72326
rect 9109 72304 9417 72324
rect 10140 72072 10192 72078
rect 10140 72014 10192 72020
rect 8392 72004 8444 72010
rect 8392 71946 8444 71952
rect 9956 71936 10008 71942
rect 9956 71878 10008 71884
rect 9968 71670 9996 71878
rect 9956 71664 10008 71670
rect 10152 71641 10180 72014
rect 9956 71606 10008 71612
rect 10138 71632 10194 71641
rect 10138 71567 10194 71576
rect 9109 71292 9417 71312
rect 9109 71290 9115 71292
rect 9171 71290 9195 71292
rect 9251 71290 9275 71292
rect 9331 71290 9355 71292
rect 9411 71290 9417 71292
rect 9171 71238 9173 71290
rect 9353 71238 9355 71290
rect 9109 71236 9115 71238
rect 9171 71236 9195 71238
rect 9251 71236 9275 71238
rect 9331 71236 9355 71238
rect 9411 71236 9417 71238
rect 9109 71216 9417 71236
rect 10140 70984 10192 70990
rect 10140 70926 10192 70932
rect 9864 70916 9916 70922
rect 9864 70858 9916 70864
rect 9109 70204 9417 70224
rect 9109 70202 9115 70204
rect 9171 70202 9195 70204
rect 9251 70202 9275 70204
rect 9331 70202 9355 70204
rect 9411 70202 9417 70204
rect 9171 70150 9173 70202
rect 9353 70150 9355 70202
rect 9109 70148 9115 70150
rect 9171 70148 9195 70150
rect 9251 70148 9275 70150
rect 9331 70148 9355 70150
rect 9411 70148 9417 70150
rect 9109 70128 9417 70148
rect 9876 70106 9904 70858
rect 9956 70848 10008 70854
rect 9956 70790 10008 70796
rect 9968 70582 9996 70790
rect 9956 70576 10008 70582
rect 10152 70553 10180 70926
rect 9956 70518 10008 70524
rect 10138 70544 10194 70553
rect 10138 70479 10194 70488
rect 9864 70100 9916 70106
rect 9864 70042 9916 70048
rect 10140 69896 10192 69902
rect 10140 69838 10192 69844
rect 10152 69465 10180 69838
rect 10138 69456 10194 69465
rect 10138 69391 10194 69400
rect 9109 69116 9417 69136
rect 9109 69114 9115 69116
rect 9171 69114 9195 69116
rect 9251 69114 9275 69116
rect 9331 69114 9355 69116
rect 9411 69114 9417 69116
rect 9171 69062 9173 69114
rect 9353 69062 9355 69114
rect 9109 69060 9115 69062
rect 9171 69060 9195 69062
rect 9251 69060 9275 69062
rect 9331 69060 9355 69062
rect 9411 69060 9417 69062
rect 9109 69040 9417 69060
rect 10140 68808 10192 68814
rect 10140 68750 10192 68756
rect 10152 68377 10180 68750
rect 10138 68368 10194 68377
rect 10138 68303 10194 68312
rect 9956 68196 10008 68202
rect 9956 68138 10008 68144
rect 8392 68128 8444 68134
rect 8392 68070 8444 68076
rect 8300 46912 8352 46918
rect 8300 46854 8352 46860
rect 8404 42702 8432 68070
rect 9109 68028 9417 68048
rect 9109 68026 9115 68028
rect 9171 68026 9195 68028
rect 9251 68026 9275 68028
rect 9331 68026 9355 68028
rect 9411 68026 9417 68028
rect 9171 67974 9173 68026
rect 9353 67974 9355 68026
rect 9109 67972 9115 67974
rect 9171 67972 9195 67974
rect 9251 67972 9275 67974
rect 9331 67972 9355 67974
rect 9411 67972 9417 67974
rect 9109 67952 9417 67972
rect 9109 66940 9417 66960
rect 9109 66938 9115 66940
rect 9171 66938 9195 66940
rect 9251 66938 9275 66940
rect 9331 66938 9355 66940
rect 9411 66938 9417 66940
rect 9171 66886 9173 66938
rect 9353 66886 9355 66938
rect 9109 66884 9115 66886
rect 9171 66884 9195 66886
rect 9251 66884 9275 66886
rect 9331 66884 9355 66886
rect 9411 66884 9417 66886
rect 9109 66864 9417 66884
rect 9968 66298 9996 68138
rect 10140 67584 10192 67590
rect 10140 67526 10192 67532
rect 10152 67289 10180 67526
rect 10138 67280 10194 67289
rect 10138 67215 10194 67224
rect 9956 66292 10008 66298
rect 9956 66234 10008 66240
rect 10140 66156 10192 66162
rect 10140 66098 10192 66104
rect 10152 66065 10180 66098
rect 10138 66056 10194 66065
rect 8484 66020 8536 66026
rect 10138 65991 10194 66000
rect 8484 65962 8536 65968
rect 8496 43246 8524 65962
rect 9109 65852 9417 65872
rect 9109 65850 9115 65852
rect 9171 65850 9195 65852
rect 9251 65850 9275 65852
rect 9331 65850 9355 65852
rect 9411 65850 9417 65852
rect 9171 65798 9173 65850
rect 9353 65798 9355 65850
rect 9109 65796 9115 65798
rect 9171 65796 9195 65798
rect 9251 65796 9275 65798
rect 9331 65796 9355 65798
rect 9411 65796 9417 65798
rect 9109 65776 9417 65796
rect 10140 65068 10192 65074
rect 10140 65010 10192 65016
rect 10152 64977 10180 65010
rect 10138 64968 10194 64977
rect 10138 64903 10194 64912
rect 9956 64864 10008 64870
rect 9956 64806 10008 64812
rect 9109 64764 9417 64784
rect 9109 64762 9115 64764
rect 9171 64762 9195 64764
rect 9251 64762 9275 64764
rect 9331 64762 9355 64764
rect 9411 64762 9417 64764
rect 9171 64710 9173 64762
rect 9353 64710 9355 64762
rect 9109 64708 9115 64710
rect 9171 64708 9195 64710
rect 9251 64708 9275 64710
rect 9331 64708 9355 64710
rect 9411 64708 9417 64710
rect 9109 64688 9417 64708
rect 9968 64394 9996 64806
rect 9956 64388 10008 64394
rect 9956 64330 10008 64336
rect 10140 63980 10192 63986
rect 10140 63922 10192 63928
rect 10152 63889 10180 63922
rect 10138 63880 10194 63889
rect 10138 63815 10194 63824
rect 9109 63676 9417 63696
rect 9109 63674 9115 63676
rect 9171 63674 9195 63676
rect 9251 63674 9275 63676
rect 9331 63674 9355 63676
rect 9411 63674 9417 63676
rect 9171 63622 9173 63674
rect 9353 63622 9355 63674
rect 9109 63620 9115 63622
rect 9171 63620 9195 63622
rect 9251 63620 9275 63622
rect 9331 63620 9355 63622
rect 9411 63620 9417 63622
rect 9109 63600 9417 63620
rect 10140 62892 10192 62898
rect 10140 62834 10192 62840
rect 10152 62801 10180 62834
rect 10138 62792 10194 62801
rect 10138 62727 10194 62736
rect 8576 62688 8628 62694
rect 8576 62630 8628 62636
rect 8484 43240 8536 43246
rect 8484 43182 8536 43188
rect 8392 42696 8444 42702
rect 8392 42638 8444 42644
rect 8588 41274 8616 62630
rect 9109 62588 9417 62608
rect 9109 62586 9115 62588
rect 9171 62586 9195 62588
rect 9251 62586 9275 62588
rect 9331 62586 9355 62588
rect 9411 62586 9417 62588
rect 9171 62534 9173 62586
rect 9353 62534 9355 62586
rect 9109 62532 9115 62534
rect 9171 62532 9195 62534
rect 9251 62532 9275 62534
rect 9331 62532 9355 62534
rect 9411 62532 9417 62534
rect 9109 62512 9417 62532
rect 9956 62212 10008 62218
rect 9956 62154 10008 62160
rect 8668 61600 8720 61606
rect 8668 61542 8720 61548
rect 8576 41268 8628 41274
rect 8576 41210 8628 41216
rect 8680 40526 8708 61542
rect 9109 61500 9417 61520
rect 9109 61498 9115 61500
rect 9171 61498 9195 61500
rect 9251 61498 9275 61500
rect 9331 61498 9355 61500
rect 9411 61498 9417 61500
rect 9171 61446 9173 61498
rect 9353 61446 9355 61498
rect 9109 61444 9115 61446
rect 9171 61444 9195 61446
rect 9251 61444 9275 61446
rect 9331 61444 9355 61446
rect 9411 61444 9417 61446
rect 9109 61424 9417 61444
rect 9968 60858 9996 62154
rect 10140 61804 10192 61810
rect 10140 61746 10192 61752
rect 10152 61713 10180 61746
rect 10138 61704 10194 61713
rect 10138 61639 10194 61648
rect 9956 60852 10008 60858
rect 9956 60794 10008 60800
rect 10140 60716 10192 60722
rect 10140 60658 10192 60664
rect 10152 60625 10180 60658
rect 10138 60616 10194 60625
rect 10138 60551 10194 60560
rect 9109 60412 9417 60432
rect 9109 60410 9115 60412
rect 9171 60410 9195 60412
rect 9251 60410 9275 60412
rect 9331 60410 9355 60412
rect 9411 60410 9417 60412
rect 9171 60358 9173 60410
rect 9353 60358 9355 60410
rect 9109 60356 9115 60358
rect 9171 60356 9195 60358
rect 9251 60356 9275 60358
rect 9331 60356 9355 60358
rect 9411 60356 9417 60358
rect 9109 60336 9417 60356
rect 10140 59628 10192 59634
rect 10140 59570 10192 59576
rect 9956 59424 10008 59430
rect 10152 59401 10180 59570
rect 9956 59366 10008 59372
rect 10138 59392 10194 59401
rect 9109 59324 9417 59344
rect 9109 59322 9115 59324
rect 9171 59322 9195 59324
rect 9251 59322 9275 59324
rect 9331 59322 9355 59324
rect 9411 59322 9417 59324
rect 9171 59270 9173 59322
rect 9353 59270 9355 59322
rect 9109 59268 9115 59270
rect 9171 59268 9195 59270
rect 9251 59268 9275 59270
rect 9331 59268 9355 59270
rect 9411 59268 9417 59270
rect 9109 59248 9417 59268
rect 9968 58954 9996 59366
rect 10138 59327 10194 59336
rect 9956 58948 10008 58954
rect 9956 58890 10008 58896
rect 10140 58540 10192 58546
rect 10140 58482 10192 58488
rect 10152 58313 10180 58482
rect 10138 58304 10194 58313
rect 9109 58236 9417 58256
rect 10138 58239 10194 58248
rect 9109 58234 9115 58236
rect 9171 58234 9195 58236
rect 9251 58234 9275 58236
rect 9331 58234 9355 58236
rect 9411 58234 9417 58236
rect 9171 58182 9173 58234
rect 9353 58182 9355 58234
rect 9109 58180 9115 58182
rect 9171 58180 9195 58182
rect 9251 58180 9275 58182
rect 9331 58180 9355 58182
rect 9411 58180 9417 58182
rect 9109 58160 9417 58180
rect 9864 57520 9916 57526
rect 9864 57462 9916 57468
rect 9109 57148 9417 57168
rect 9109 57146 9115 57148
rect 9171 57146 9195 57148
rect 9251 57146 9275 57148
rect 9331 57146 9355 57148
rect 9411 57146 9417 57148
rect 9171 57094 9173 57146
rect 9353 57094 9355 57146
rect 9109 57092 9115 57094
rect 9171 57092 9195 57094
rect 9251 57092 9275 57094
rect 9331 57092 9355 57094
rect 9411 57092 9417 57094
rect 9109 57072 9417 57092
rect 9109 56060 9417 56080
rect 9109 56058 9115 56060
rect 9171 56058 9195 56060
rect 9251 56058 9275 56060
rect 9331 56058 9355 56060
rect 9411 56058 9417 56060
rect 9171 56006 9173 56058
rect 9353 56006 9355 56058
rect 9109 56004 9115 56006
rect 9171 56004 9195 56006
rect 9251 56004 9275 56006
rect 9331 56004 9355 56006
rect 9411 56004 9417 56006
rect 9109 55984 9417 56004
rect 9876 55418 9904 57462
rect 10140 57452 10192 57458
rect 10140 57394 10192 57400
rect 9956 57248 10008 57254
rect 10152 57225 10180 57394
rect 9956 57190 10008 57196
rect 10138 57216 10194 57225
rect 9968 57050 9996 57190
rect 10138 57151 10194 57160
rect 9956 57044 10008 57050
rect 9956 56986 10008 56992
rect 9956 56772 10008 56778
rect 9956 56714 10008 56720
rect 9968 56506 9996 56714
rect 9956 56500 10008 56506
rect 9956 56442 10008 56448
rect 10140 56364 10192 56370
rect 10140 56306 10192 56312
rect 10152 56137 10180 56306
rect 10138 56128 10194 56137
rect 10138 56063 10194 56072
rect 9864 55412 9916 55418
rect 9864 55354 9916 55360
rect 10140 55276 10192 55282
rect 10140 55218 10192 55224
rect 10152 55049 10180 55218
rect 10138 55040 10194 55049
rect 9109 54972 9417 54992
rect 10138 54975 10194 54984
rect 9109 54970 9115 54972
rect 9171 54970 9195 54972
rect 9251 54970 9275 54972
rect 9331 54970 9355 54972
rect 9411 54970 9417 54972
rect 9171 54918 9173 54970
rect 9353 54918 9355 54970
rect 9109 54916 9115 54918
rect 9171 54916 9195 54918
rect 9251 54916 9275 54918
rect 9331 54916 9355 54918
rect 9411 54916 9417 54918
rect 9109 54896 9417 54916
rect 10140 54188 10192 54194
rect 10140 54130 10192 54136
rect 9956 53984 10008 53990
rect 10152 53961 10180 54130
rect 9956 53926 10008 53932
rect 10138 53952 10194 53961
rect 9109 53884 9417 53904
rect 9109 53882 9115 53884
rect 9171 53882 9195 53884
rect 9251 53882 9275 53884
rect 9331 53882 9355 53884
rect 9411 53882 9417 53884
rect 9171 53830 9173 53882
rect 9353 53830 9355 53882
rect 9109 53828 9115 53830
rect 9171 53828 9195 53830
rect 9251 53828 9275 53830
rect 9331 53828 9355 53830
rect 9411 53828 9417 53830
rect 9109 53808 9417 53828
rect 9968 53174 9996 53926
rect 10138 53887 10194 53896
rect 9956 53168 10008 53174
rect 9956 53110 10008 53116
rect 10140 53100 10192 53106
rect 10140 53042 10192 53048
rect 9956 52896 10008 52902
rect 9956 52838 10008 52844
rect 9109 52796 9417 52816
rect 9109 52794 9115 52796
rect 9171 52794 9195 52796
rect 9251 52794 9275 52796
rect 9331 52794 9355 52796
rect 9411 52794 9417 52796
rect 9171 52742 9173 52794
rect 9353 52742 9355 52794
rect 9109 52740 9115 52742
rect 9171 52740 9195 52742
rect 9251 52740 9275 52742
rect 9331 52740 9355 52742
rect 9411 52740 9417 52742
rect 9109 52720 9417 52740
rect 9968 52562 9996 52838
rect 10152 52737 10180 53042
rect 10138 52728 10194 52737
rect 10138 52663 10194 52672
rect 9956 52556 10008 52562
rect 9956 52498 10008 52504
rect 10140 52012 10192 52018
rect 10140 51954 10192 51960
rect 9956 51808 10008 51814
rect 9956 51750 10008 51756
rect 9109 51708 9417 51728
rect 9109 51706 9115 51708
rect 9171 51706 9195 51708
rect 9251 51706 9275 51708
rect 9331 51706 9355 51708
rect 9411 51706 9417 51708
rect 9171 51654 9173 51706
rect 9353 51654 9355 51706
rect 9109 51652 9115 51654
rect 9171 51652 9195 51654
rect 9251 51652 9275 51654
rect 9331 51652 9355 51654
rect 9411 51652 9417 51654
rect 9109 51632 9417 51652
rect 9864 51604 9916 51610
rect 9864 51546 9916 51552
rect 9876 51066 9904 51546
rect 9968 51338 9996 51750
rect 10152 51649 10180 51954
rect 10138 51640 10194 51649
rect 10138 51575 10194 51584
rect 9956 51332 10008 51338
rect 9956 51274 10008 51280
rect 9864 51060 9916 51066
rect 9864 51002 9916 51008
rect 10140 50924 10192 50930
rect 10140 50866 10192 50872
rect 9109 50620 9417 50640
rect 9109 50618 9115 50620
rect 9171 50618 9195 50620
rect 9251 50618 9275 50620
rect 9331 50618 9355 50620
rect 9411 50618 9417 50620
rect 9171 50566 9173 50618
rect 9353 50566 9355 50618
rect 9109 50564 9115 50566
rect 9171 50564 9195 50566
rect 9251 50564 9275 50566
rect 9331 50564 9355 50566
rect 9411 50564 9417 50566
rect 9109 50544 9417 50564
rect 10152 50561 10180 50866
rect 10138 50552 10194 50561
rect 10138 50487 10194 50496
rect 9956 50244 10008 50250
rect 9956 50186 10008 50192
rect 9968 49978 9996 50186
rect 9956 49972 10008 49978
rect 9956 49914 10008 49920
rect 10140 49700 10192 49706
rect 10140 49642 10192 49648
rect 9109 49532 9417 49552
rect 9109 49530 9115 49532
rect 9171 49530 9195 49532
rect 9251 49530 9275 49532
rect 9331 49530 9355 49532
rect 9411 49530 9417 49532
rect 9171 49478 9173 49530
rect 9353 49478 9355 49530
rect 9109 49476 9115 49478
rect 9171 49476 9195 49478
rect 9251 49476 9275 49478
rect 9331 49476 9355 49478
rect 9411 49476 9417 49478
rect 9109 49456 9417 49476
rect 10152 49473 10180 49642
rect 10138 49464 10194 49473
rect 10138 49399 10194 49408
rect 10140 48748 10192 48754
rect 10140 48690 10192 48696
rect 9109 48444 9417 48464
rect 9109 48442 9115 48444
rect 9171 48442 9195 48444
rect 9251 48442 9275 48444
rect 9331 48442 9355 48444
rect 9411 48442 9417 48444
rect 9171 48390 9173 48442
rect 9353 48390 9355 48442
rect 9109 48388 9115 48390
rect 9171 48388 9195 48390
rect 9251 48388 9275 48390
rect 9331 48388 9355 48390
rect 9411 48388 9417 48390
rect 9109 48368 9417 48388
rect 10152 48385 10180 48690
rect 10138 48376 10194 48385
rect 10138 48311 10194 48320
rect 10140 47660 10192 47666
rect 10140 47602 10192 47608
rect 9109 47356 9417 47376
rect 9109 47354 9115 47356
rect 9171 47354 9195 47356
rect 9251 47354 9275 47356
rect 9331 47354 9355 47356
rect 9411 47354 9417 47356
rect 9171 47302 9173 47354
rect 9353 47302 9355 47354
rect 9109 47300 9115 47302
rect 9171 47300 9195 47302
rect 9251 47300 9275 47302
rect 9331 47300 9355 47302
rect 9411 47300 9417 47302
rect 9109 47280 9417 47300
rect 10152 47297 10180 47602
rect 10138 47288 10194 47297
rect 10138 47223 10194 47232
rect 10140 46572 10192 46578
rect 10140 46514 10192 46520
rect 9956 46368 10008 46374
rect 9956 46310 10008 46316
rect 9109 46268 9417 46288
rect 9109 46266 9115 46268
rect 9171 46266 9195 46268
rect 9251 46266 9275 46268
rect 9331 46266 9355 46268
rect 9411 46266 9417 46268
rect 9171 46214 9173 46266
rect 9353 46214 9355 46266
rect 9109 46212 9115 46214
rect 9171 46212 9195 46214
rect 9251 46212 9275 46214
rect 9331 46212 9355 46214
rect 9411 46212 9417 46214
rect 9109 46192 9417 46212
rect 9864 45280 9916 45286
rect 9864 45222 9916 45228
rect 9109 45180 9417 45200
rect 9109 45178 9115 45180
rect 9171 45178 9195 45180
rect 9251 45178 9275 45180
rect 9331 45178 9355 45180
rect 9411 45178 9417 45180
rect 9171 45126 9173 45178
rect 9353 45126 9355 45178
rect 9109 45124 9115 45126
rect 9171 45124 9195 45126
rect 9251 45124 9275 45126
rect 9331 45124 9355 45126
rect 9411 45124 9417 45126
rect 9109 45104 9417 45124
rect 9109 44092 9417 44112
rect 9109 44090 9115 44092
rect 9171 44090 9195 44092
rect 9251 44090 9275 44092
rect 9331 44090 9355 44092
rect 9411 44090 9417 44092
rect 9171 44038 9173 44090
rect 9353 44038 9355 44090
rect 9109 44036 9115 44038
rect 9171 44036 9195 44038
rect 9251 44036 9275 44038
rect 9331 44036 9355 44038
rect 9411 44036 9417 44038
rect 9109 44016 9417 44036
rect 9876 43450 9904 45222
rect 9968 44470 9996 46310
rect 10152 46073 10180 46514
rect 10138 46064 10194 46073
rect 10138 45999 10194 46008
rect 10140 45484 10192 45490
rect 10140 45426 10192 45432
rect 10152 44985 10180 45426
rect 10138 44976 10194 44985
rect 10138 44911 10194 44920
rect 9956 44464 10008 44470
rect 9956 44406 10008 44412
rect 10140 44396 10192 44402
rect 10140 44338 10192 44344
rect 9956 44192 10008 44198
rect 9956 44134 10008 44140
rect 9968 43722 9996 44134
rect 10152 43897 10180 44338
rect 10138 43888 10194 43897
rect 10138 43823 10194 43832
rect 9956 43716 10008 43722
rect 9956 43658 10008 43664
rect 9864 43444 9916 43450
rect 9864 43386 9916 43392
rect 9864 43308 9916 43314
rect 9864 43250 9916 43256
rect 9109 43004 9417 43024
rect 9109 43002 9115 43004
rect 9171 43002 9195 43004
rect 9251 43002 9275 43004
rect 9331 43002 9355 43004
rect 9411 43002 9417 43004
rect 9171 42950 9173 43002
rect 9353 42950 9355 43002
rect 9109 42948 9115 42950
rect 9171 42948 9195 42950
rect 9251 42948 9275 42950
rect 9331 42948 9355 42950
rect 9411 42948 9417 42950
rect 9109 42928 9417 42948
rect 9876 42770 9904 43250
rect 10048 43104 10100 43110
rect 10048 43046 10100 43052
rect 10060 42809 10088 43046
rect 10046 42800 10102 42809
rect 9864 42764 9916 42770
rect 10046 42735 10102 42744
rect 9864 42706 9916 42712
rect 10048 42016 10100 42022
rect 10048 41958 10100 41964
rect 9109 41916 9417 41936
rect 9109 41914 9115 41916
rect 9171 41914 9195 41916
rect 9251 41914 9275 41916
rect 9331 41914 9355 41916
rect 9411 41914 9417 41916
rect 9171 41862 9173 41914
rect 9353 41862 9355 41914
rect 9109 41860 9115 41862
rect 9171 41860 9195 41862
rect 9251 41860 9275 41862
rect 9331 41860 9355 41862
rect 9411 41860 9417 41862
rect 9109 41840 9417 41860
rect 10060 41721 10088 41958
rect 10046 41712 10102 41721
rect 10046 41647 10102 41656
rect 10048 40928 10100 40934
rect 10048 40870 10100 40876
rect 9109 40828 9417 40848
rect 9109 40826 9115 40828
rect 9171 40826 9195 40828
rect 9251 40826 9275 40828
rect 9331 40826 9355 40828
rect 9411 40826 9417 40828
rect 9171 40774 9173 40826
rect 9353 40774 9355 40826
rect 9109 40772 9115 40774
rect 9171 40772 9195 40774
rect 9251 40772 9275 40774
rect 9331 40772 9355 40774
rect 9411 40772 9417 40774
rect 9109 40752 9417 40772
rect 10060 40633 10088 40870
rect 10046 40624 10102 40633
rect 10046 40559 10102 40568
rect 8668 40520 8720 40526
rect 8668 40462 8720 40468
rect 9109 39740 9417 39760
rect 9109 39738 9115 39740
rect 9171 39738 9195 39740
rect 9251 39738 9275 39740
rect 9331 39738 9355 39740
rect 9411 39738 9417 39740
rect 9171 39686 9173 39738
rect 9353 39686 9355 39738
rect 9109 39684 9115 39686
rect 9171 39684 9195 39686
rect 9251 39684 9275 39686
rect 9331 39684 9355 39686
rect 9411 39684 9417 39686
rect 9109 39664 9417 39684
rect 9864 39432 9916 39438
rect 9864 39374 9916 39380
rect 10046 39400 10102 39409
rect 9876 38758 9904 39374
rect 10046 39335 10102 39344
rect 10060 39302 10088 39335
rect 10048 39296 10100 39302
rect 10048 39238 10100 39244
rect 9864 38752 9916 38758
rect 9864 38694 9916 38700
rect 9109 38652 9417 38672
rect 9109 38650 9115 38652
rect 9171 38650 9195 38652
rect 9251 38650 9275 38652
rect 9331 38650 9355 38652
rect 9411 38650 9417 38652
rect 9171 38598 9173 38650
rect 9353 38598 9355 38650
rect 9109 38596 9115 38598
rect 9171 38596 9195 38598
rect 9251 38596 9275 38598
rect 9331 38596 9355 38598
rect 9411 38596 9417 38598
rect 9109 38576 9417 38596
rect 10046 38312 10102 38321
rect 10046 38247 10102 38256
rect 10060 38214 10088 38247
rect 10048 38208 10100 38214
rect 10048 38150 10100 38156
rect 9864 37664 9916 37670
rect 9864 37606 9916 37612
rect 9109 37564 9417 37584
rect 9109 37562 9115 37564
rect 9171 37562 9195 37564
rect 9251 37562 9275 37564
rect 9331 37562 9355 37564
rect 9411 37562 9417 37564
rect 9171 37510 9173 37562
rect 9353 37510 9355 37562
rect 9109 37508 9115 37510
rect 9171 37508 9195 37510
rect 9251 37508 9275 37510
rect 9331 37508 9355 37510
rect 9411 37508 9417 37510
rect 9109 37488 9417 37508
rect 9876 37262 9904 37606
rect 9864 37256 9916 37262
rect 9864 37198 9916 37204
rect 10046 37224 10102 37233
rect 10046 37159 10102 37168
rect 10060 37126 10088 37159
rect 10048 37120 10100 37126
rect 10048 37062 10100 37068
rect 9864 36576 9916 36582
rect 9864 36518 9916 36524
rect 9109 36476 9417 36496
rect 9109 36474 9115 36476
rect 9171 36474 9195 36476
rect 9251 36474 9275 36476
rect 9331 36474 9355 36476
rect 9411 36474 9417 36476
rect 9171 36422 9173 36474
rect 9353 36422 9355 36474
rect 9109 36420 9115 36422
rect 9171 36420 9195 36422
rect 9251 36420 9275 36422
rect 9331 36420 9355 36422
rect 9411 36420 9417 36422
rect 9109 36400 9417 36420
rect 9876 36174 9904 36518
rect 9864 36168 9916 36174
rect 9864 36110 9916 36116
rect 10046 36136 10102 36145
rect 10046 36071 10102 36080
rect 10060 36038 10088 36071
rect 9864 36032 9916 36038
rect 9864 35974 9916 35980
rect 10048 36032 10100 36038
rect 10048 35974 10100 35980
rect 9109 35388 9417 35408
rect 9109 35386 9115 35388
rect 9171 35386 9195 35388
rect 9251 35386 9275 35388
rect 9331 35386 9355 35388
rect 9411 35386 9417 35388
rect 9171 35334 9173 35386
rect 9353 35334 9355 35386
rect 9109 35332 9115 35334
rect 9171 35332 9195 35334
rect 9251 35332 9275 35334
rect 9331 35332 9355 35334
rect 9411 35332 9417 35334
rect 9109 35312 9417 35332
rect 9876 35086 9904 35974
rect 9864 35080 9916 35086
rect 9864 35022 9916 35028
rect 10046 35048 10102 35057
rect 10046 34983 10102 34992
rect 10060 34950 10088 34983
rect 10048 34944 10100 34950
rect 10048 34886 10100 34892
rect 9109 34300 9417 34320
rect 9109 34298 9115 34300
rect 9171 34298 9195 34300
rect 9251 34298 9275 34300
rect 9331 34298 9355 34300
rect 9411 34298 9417 34300
rect 9171 34246 9173 34298
rect 9353 34246 9355 34298
rect 9109 34244 9115 34246
rect 9171 34244 9195 34246
rect 9251 34244 9275 34246
rect 9331 34244 9355 34246
rect 9411 34244 9417 34246
rect 9109 34224 9417 34244
rect 9864 33992 9916 33998
rect 9864 33934 9916 33940
rect 10046 33960 10102 33969
rect 9876 33318 9904 33934
rect 10046 33895 10102 33904
rect 10060 33862 10088 33895
rect 10048 33856 10100 33862
rect 10048 33798 10100 33804
rect 9864 33312 9916 33318
rect 9864 33254 9916 33260
rect 9109 33212 9417 33232
rect 9109 33210 9115 33212
rect 9171 33210 9195 33212
rect 9251 33210 9275 33212
rect 9331 33210 9355 33212
rect 9411 33210 9417 33212
rect 9171 33158 9173 33210
rect 9353 33158 9355 33210
rect 9109 33156 9115 33158
rect 9171 33156 9195 33158
rect 9251 33156 9275 33158
rect 9331 33156 9355 33158
rect 9411 33156 9417 33158
rect 9109 33136 9417 33156
rect 10048 32768 10100 32774
rect 10046 32736 10048 32745
rect 10100 32736 10102 32745
rect 10046 32671 10102 32680
rect 9109 32124 9417 32144
rect 9109 32122 9115 32124
rect 9171 32122 9195 32124
rect 9251 32122 9275 32124
rect 9331 32122 9355 32124
rect 9411 32122 9417 32124
rect 9171 32070 9173 32122
rect 9353 32070 9355 32122
rect 9109 32068 9115 32070
rect 9171 32068 9195 32070
rect 9251 32068 9275 32070
rect 9331 32068 9355 32070
rect 9411 32068 9417 32070
rect 9109 32048 9417 32068
rect 10048 31680 10100 31686
rect 10046 31648 10048 31657
rect 10100 31648 10102 31657
rect 10046 31583 10102 31592
rect 9864 31136 9916 31142
rect 9864 31078 9916 31084
rect 9109 31036 9417 31056
rect 9109 31034 9115 31036
rect 9171 31034 9195 31036
rect 9251 31034 9275 31036
rect 9331 31034 9355 31036
rect 9411 31034 9417 31036
rect 9171 30982 9173 31034
rect 9353 30982 9355 31034
rect 9109 30980 9115 30982
rect 9171 30980 9195 30982
rect 9251 30980 9275 30982
rect 9331 30980 9355 30982
rect 9411 30980 9417 30982
rect 9109 30960 9417 30980
rect 9876 30734 9904 31078
rect 9864 30728 9916 30734
rect 9864 30670 9916 30676
rect 9864 30592 9916 30598
rect 10048 30592 10100 30598
rect 9864 30534 9916 30540
rect 10046 30560 10048 30569
rect 10100 30560 10102 30569
rect 9109 29948 9417 29968
rect 9109 29946 9115 29948
rect 9171 29946 9195 29948
rect 9251 29946 9275 29948
rect 9331 29946 9355 29948
rect 9411 29946 9417 29948
rect 9171 29894 9173 29946
rect 9353 29894 9355 29946
rect 9109 29892 9115 29894
rect 9171 29892 9195 29894
rect 9251 29892 9275 29894
rect 9331 29892 9355 29894
rect 9411 29892 9417 29894
rect 9109 29872 9417 29892
rect 9876 29646 9904 30534
rect 10046 30495 10102 30504
rect 9864 29640 9916 29646
rect 9864 29582 9916 29588
rect 10048 29504 10100 29510
rect 10046 29472 10048 29481
rect 10100 29472 10102 29481
rect 10046 29407 10102 29416
rect 9109 28860 9417 28880
rect 9109 28858 9115 28860
rect 9171 28858 9195 28860
rect 9251 28858 9275 28860
rect 9331 28858 9355 28860
rect 9411 28858 9417 28860
rect 9171 28806 9173 28858
rect 9353 28806 9355 28858
rect 9109 28804 9115 28806
rect 9171 28804 9195 28806
rect 9251 28804 9275 28806
rect 9331 28804 9355 28806
rect 9411 28804 9417 28806
rect 9109 28784 9417 28804
rect 10048 28416 10100 28422
rect 10046 28384 10048 28393
rect 10100 28384 10102 28393
rect 10046 28319 10102 28328
rect 9109 27772 9417 27792
rect 9109 27770 9115 27772
rect 9171 27770 9195 27772
rect 9251 27770 9275 27772
rect 9331 27770 9355 27772
rect 9411 27770 9417 27772
rect 9171 27718 9173 27770
rect 9353 27718 9355 27770
rect 9109 27716 9115 27718
rect 9171 27716 9195 27718
rect 9251 27716 9275 27718
rect 9331 27716 9355 27718
rect 9411 27716 9417 27718
rect 9109 27696 9417 27716
rect 10048 27328 10100 27334
rect 10046 27296 10048 27305
rect 10100 27296 10102 27305
rect 10046 27231 10102 27240
rect 9864 26784 9916 26790
rect 9864 26726 9916 26732
rect 9109 26684 9417 26704
rect 9109 26682 9115 26684
rect 9171 26682 9195 26684
rect 9251 26682 9275 26684
rect 9331 26682 9355 26684
rect 9411 26682 9417 26684
rect 9171 26630 9173 26682
rect 9353 26630 9355 26682
rect 9109 26628 9115 26630
rect 9171 26628 9195 26630
rect 9251 26628 9275 26630
rect 9331 26628 9355 26630
rect 9411 26628 9417 26630
rect 9109 26608 9417 26628
rect 9876 26382 9904 26726
rect 9956 26512 10008 26518
rect 9956 26454 10008 26460
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 9109 25596 9417 25616
rect 9109 25594 9115 25596
rect 9171 25594 9195 25596
rect 9251 25594 9275 25596
rect 9331 25594 9355 25596
rect 9411 25594 9417 25596
rect 9171 25542 9173 25594
rect 9353 25542 9355 25594
rect 9109 25540 9115 25542
rect 9171 25540 9195 25542
rect 9251 25540 9275 25542
rect 9331 25540 9355 25542
rect 9411 25540 9417 25542
rect 9109 25520 9417 25540
rect 9109 24508 9417 24528
rect 9109 24506 9115 24508
rect 9171 24506 9195 24508
rect 9251 24506 9275 24508
rect 9331 24506 9355 24508
rect 9411 24506 9417 24508
rect 9171 24454 9173 24506
rect 9353 24454 9355 24506
rect 9109 24452 9115 24454
rect 9171 24452 9195 24454
rect 9251 24452 9275 24454
rect 9331 24452 9355 24454
rect 9411 24452 9417 24454
rect 9109 24432 9417 24452
rect 9784 24206 9812 26250
rect 9968 25294 9996 26454
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 10060 26081 10088 26182
rect 10046 26072 10102 26081
rect 10046 26007 10102 26016
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 10060 24993 10088 25094
rect 10046 24984 10102 24993
rect 10046 24919 10102 24928
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 10060 23905 10088 24006
rect 10046 23896 10102 23905
rect 10046 23831 10102 23840
rect 9109 23420 9417 23440
rect 9109 23418 9115 23420
rect 9171 23418 9195 23420
rect 9251 23418 9275 23420
rect 9331 23418 9355 23420
rect 9411 23418 9417 23420
rect 9171 23366 9173 23418
rect 9353 23366 9355 23418
rect 9109 23364 9115 23366
rect 9171 23364 9195 23366
rect 9251 23364 9275 23366
rect 9331 23364 9355 23366
rect 9411 23364 9417 23366
rect 9109 23344 9417 23364
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 10060 22817 10088 22918
rect 10046 22808 10102 22817
rect 9864 22772 9916 22778
rect 10046 22743 10102 22752
rect 9864 22714 9916 22720
rect 9109 22332 9417 22352
rect 9109 22330 9115 22332
rect 9171 22330 9195 22332
rect 9251 22330 9275 22332
rect 9331 22330 9355 22332
rect 9411 22330 9417 22332
rect 9171 22278 9173 22330
rect 9353 22278 9355 22330
rect 9109 22276 9115 22278
rect 9171 22276 9195 22278
rect 9251 22276 9275 22278
rect 9331 22276 9355 22278
rect 9411 22276 9417 22278
rect 9109 22256 9417 22276
rect 9876 22030 9904 22714
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 9109 21244 9417 21264
rect 9109 21242 9115 21244
rect 9171 21242 9195 21244
rect 9251 21242 9275 21244
rect 9331 21242 9355 21244
rect 9411 21242 9417 21244
rect 9171 21190 9173 21242
rect 9353 21190 9355 21242
rect 9109 21188 9115 21190
rect 9171 21188 9195 21190
rect 9251 21188 9275 21190
rect 9331 21188 9355 21190
rect 9411 21188 9417 21190
rect 9109 21168 9417 21188
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9109 20156 9417 20176
rect 9109 20154 9115 20156
rect 9171 20154 9195 20156
rect 9251 20154 9275 20156
rect 9331 20154 9355 20156
rect 9411 20154 9417 20156
rect 9171 20102 9173 20154
rect 9353 20102 9355 20154
rect 9109 20100 9115 20102
rect 9171 20100 9195 20102
rect 9251 20100 9275 20102
rect 9331 20100 9355 20102
rect 9411 20100 9417 20102
rect 9109 20080 9417 20100
rect 9784 19854 9812 21082
rect 9876 20942 9904 21830
rect 10060 21729 10088 21830
rect 10046 21720 10102 21729
rect 10046 21655 10102 21664
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 10060 20641 10088 20742
rect 10046 20632 10102 20641
rect 10046 20567 10102 20576
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10060 19417 10088 19654
rect 10046 19408 10102 19417
rect 10046 19343 10102 19352
rect 9109 19068 9417 19088
rect 9109 19066 9115 19068
rect 9171 19066 9195 19068
rect 9251 19066 9275 19068
rect 9331 19066 9355 19068
rect 9411 19066 9417 19068
rect 9171 19014 9173 19066
rect 9353 19014 9355 19066
rect 9109 19012 9115 19014
rect 9171 19012 9195 19014
rect 9251 19012 9275 19014
rect 9331 19012 9355 19014
rect 9411 19012 9417 19014
rect 9109 18992 9417 19012
rect 7840 18692 7892 18698
rect 7840 18634 7892 18640
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 7477 18524 7785 18544
rect 7477 18522 7483 18524
rect 7539 18522 7563 18524
rect 7619 18522 7643 18524
rect 7699 18522 7723 18524
rect 7779 18522 7785 18524
rect 7539 18470 7541 18522
rect 7721 18470 7723 18522
rect 7477 18468 7483 18470
rect 7539 18468 7563 18470
rect 7619 18468 7643 18470
rect 7699 18468 7723 18470
rect 7779 18468 7785 18470
rect 7477 18448 7785 18468
rect 10060 18329 10088 18566
rect 10046 18320 10102 18329
rect 10046 18255 10102 18264
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9109 17980 9417 18000
rect 9109 17978 9115 17980
rect 9171 17978 9195 17980
rect 9251 17978 9275 17980
rect 9331 17978 9355 17980
rect 9411 17978 9417 17980
rect 9171 17926 9173 17978
rect 9353 17926 9355 17978
rect 9109 17924 9115 17926
rect 9171 17924 9195 17926
rect 9251 17924 9275 17926
rect 9331 17924 9355 17926
rect 9411 17924 9417 17926
rect 9109 17904 9417 17924
rect 7477 17436 7785 17456
rect 7477 17434 7483 17436
rect 7539 17434 7563 17436
rect 7619 17434 7643 17436
rect 7699 17434 7723 17436
rect 7779 17434 7785 17436
rect 7539 17382 7541 17434
rect 7721 17382 7723 17434
rect 7477 17380 7483 17382
rect 7539 17380 7563 17382
rect 7619 17380 7643 17382
rect 7699 17380 7723 17382
rect 7779 17380 7785 17382
rect 7477 17360 7785 17380
rect 9109 16892 9417 16912
rect 9109 16890 9115 16892
rect 9171 16890 9195 16892
rect 9251 16890 9275 16892
rect 9331 16890 9355 16892
rect 9411 16890 9417 16892
rect 9171 16838 9173 16890
rect 9353 16838 9355 16890
rect 9109 16836 9115 16838
rect 9171 16836 9195 16838
rect 9251 16836 9275 16838
rect 9331 16836 9355 16838
rect 9411 16836 9417 16838
rect 9109 16816 9417 16836
rect 9784 16590 9812 18090
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 17678 9904 18022
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10060 17241 10088 17478
rect 10046 17232 10102 17241
rect 10046 17167 10102 17176
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 7477 16348 7785 16368
rect 7477 16346 7483 16348
rect 7539 16346 7563 16348
rect 7619 16346 7643 16348
rect 7699 16346 7723 16348
rect 7779 16346 7785 16348
rect 7539 16294 7541 16346
rect 7721 16294 7723 16346
rect 7477 16292 7483 16294
rect 7539 16292 7563 16294
rect 7619 16292 7643 16294
rect 7699 16292 7723 16294
rect 7779 16292 7785 16294
rect 7477 16272 7785 16292
rect 9109 15804 9417 15824
rect 9109 15802 9115 15804
rect 9171 15802 9195 15804
rect 9251 15802 9275 15804
rect 9331 15802 9355 15804
rect 9411 15802 9417 15804
rect 9171 15750 9173 15802
rect 9353 15750 9355 15802
rect 9109 15748 9115 15750
rect 9171 15748 9195 15750
rect 9251 15748 9275 15750
rect 9331 15748 9355 15750
rect 9411 15748 9417 15750
rect 9109 15728 9417 15748
rect 9876 15502 9904 16934
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10060 16153 10088 16390
rect 10046 16144 10102 16153
rect 10046 16079 10102 16088
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 7477 15260 7785 15280
rect 7477 15258 7483 15260
rect 7539 15258 7563 15260
rect 7619 15258 7643 15260
rect 7699 15258 7723 15260
rect 7779 15258 7785 15260
rect 7539 15206 7541 15258
rect 7721 15206 7723 15258
rect 7477 15204 7483 15206
rect 7539 15204 7563 15206
rect 7619 15204 7643 15206
rect 7699 15204 7723 15206
rect 7779 15204 7785 15206
rect 7477 15184 7785 15204
rect 10060 15065 10088 15302
rect 10046 15056 10102 15065
rect 10046 14991 10102 15000
rect 9109 14716 9417 14736
rect 9109 14714 9115 14716
rect 9171 14714 9195 14716
rect 9251 14714 9275 14716
rect 9331 14714 9355 14716
rect 9411 14714 9417 14716
rect 9171 14662 9173 14714
rect 9353 14662 9355 14714
rect 9109 14660 9115 14662
rect 9171 14660 9195 14662
rect 9251 14660 9275 14662
rect 9331 14660 9355 14662
rect 9411 14660 9417 14662
rect 9109 14640 9417 14660
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 7477 14172 7785 14192
rect 7477 14170 7483 14172
rect 7539 14170 7563 14172
rect 7619 14170 7643 14172
rect 7699 14170 7723 14172
rect 7779 14170 7785 14172
rect 7539 14118 7541 14170
rect 7721 14118 7723 14170
rect 7477 14116 7483 14118
rect 7539 14116 7563 14118
rect 7619 14116 7643 14118
rect 7699 14116 7723 14118
rect 7779 14116 7785 14118
rect 7477 14096 7785 14116
rect 10060 13977 10088 14214
rect 10046 13968 10102 13977
rect 10046 13903 10102 13912
rect 9109 13628 9417 13648
rect 9109 13626 9115 13628
rect 9171 13626 9195 13628
rect 9251 13626 9275 13628
rect 9331 13626 9355 13628
rect 9411 13626 9417 13628
rect 9171 13574 9173 13626
rect 9353 13574 9355 13626
rect 9109 13572 9115 13574
rect 9171 13572 9195 13574
rect 9251 13572 9275 13574
rect 9331 13572 9355 13574
rect 9411 13572 9417 13574
rect 9109 13552 9417 13572
rect 7477 13084 7785 13104
rect 7477 13082 7483 13084
rect 7539 13082 7563 13084
rect 7619 13082 7643 13084
rect 7699 13082 7723 13084
rect 7779 13082 7785 13084
rect 7539 13030 7541 13082
rect 7721 13030 7723 13082
rect 7477 13028 7483 13030
rect 7539 13028 7563 13030
rect 7619 13028 7643 13030
rect 7699 13028 7723 13030
rect 7779 13028 7785 13030
rect 7477 13008 7785 13028
rect 10046 12744 10102 12753
rect 10046 12679 10048 12688
rect 10100 12679 10102 12688
rect 10048 12650 10100 12656
rect 9109 12540 9417 12560
rect 9109 12538 9115 12540
rect 9171 12538 9195 12540
rect 9251 12538 9275 12540
rect 9331 12538 9355 12540
rect 9411 12538 9417 12540
rect 9171 12486 9173 12538
rect 9353 12486 9355 12538
rect 9109 12484 9115 12486
rect 9171 12484 9195 12486
rect 9251 12484 9275 12486
rect 9331 12484 9355 12486
rect 9411 12484 9417 12486
rect 9109 12464 9417 12484
rect 7477 11996 7785 12016
rect 7477 11994 7483 11996
rect 7539 11994 7563 11996
rect 7619 11994 7643 11996
rect 7699 11994 7723 11996
rect 7779 11994 7785 11996
rect 7539 11942 7541 11994
rect 7721 11942 7723 11994
rect 7477 11940 7483 11942
rect 7539 11940 7563 11942
rect 7619 11940 7643 11942
rect 7699 11940 7723 11942
rect 7779 11940 7785 11942
rect 7477 11920 7785 11940
rect 10046 11656 10102 11665
rect 10046 11591 10048 11600
rect 10100 11591 10102 11600
rect 10048 11562 10100 11568
rect 9109 11452 9417 11472
rect 9109 11450 9115 11452
rect 9171 11450 9195 11452
rect 9251 11450 9275 11452
rect 9331 11450 9355 11452
rect 9411 11450 9417 11452
rect 9171 11398 9173 11450
rect 9353 11398 9355 11450
rect 9109 11396 9115 11398
rect 9171 11396 9195 11398
rect 9251 11396 9275 11398
rect 9331 11396 9355 11398
rect 9411 11396 9417 11398
rect 9109 11376 9417 11396
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 7477 10908 7785 10928
rect 7477 10906 7483 10908
rect 7539 10906 7563 10908
rect 7619 10906 7643 10908
rect 7699 10906 7723 10908
rect 7779 10906 7785 10908
rect 7539 10854 7541 10906
rect 7721 10854 7723 10906
rect 7477 10852 7483 10854
rect 7539 10852 7563 10854
rect 7619 10852 7643 10854
rect 7699 10852 7723 10854
rect 7779 10852 7785 10854
rect 7477 10832 7785 10852
rect 9876 10674 9904 11018
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 10046 10568 10102 10577
rect 10046 10503 10048 10512
rect 10100 10503 10102 10512
rect 10048 10474 10100 10480
rect 9109 10364 9417 10384
rect 9109 10362 9115 10364
rect 9171 10362 9195 10364
rect 9251 10362 9275 10364
rect 9331 10362 9355 10364
rect 9411 10362 9417 10364
rect 9171 10310 9173 10362
rect 9353 10310 9355 10362
rect 9109 10308 9115 10310
rect 9171 10308 9195 10310
rect 9251 10308 9275 10310
rect 9331 10308 9355 10310
rect 9411 10308 9417 10310
rect 9109 10288 9417 10308
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 7477 9820 7785 9840
rect 7477 9818 7483 9820
rect 7539 9818 7563 9820
rect 7619 9818 7643 9820
rect 7699 9818 7723 9820
rect 7779 9818 7785 9820
rect 7539 9766 7541 9818
rect 7721 9766 7723 9818
rect 7477 9764 7483 9766
rect 7539 9764 7563 9766
rect 7619 9764 7643 9766
rect 7699 9764 7723 9766
rect 7779 9764 7785 9766
rect 7477 9744 7785 9764
rect 9876 9722 9904 9862
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 10046 9480 10102 9489
rect 10046 9415 10048 9424
rect 10100 9415 10102 9424
rect 10048 9386 10100 9392
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9109 9276 9417 9296
rect 9109 9274 9115 9276
rect 9171 9274 9195 9276
rect 9251 9274 9275 9276
rect 9331 9274 9355 9276
rect 9411 9274 9417 9276
rect 9171 9222 9173 9274
rect 9353 9222 9355 9274
rect 9109 9220 9115 9222
rect 9171 9220 9195 9222
rect 9251 9220 9275 9222
rect 9331 9220 9355 9222
rect 9411 9220 9417 9222
rect 9109 9200 9417 9220
rect 7477 8732 7785 8752
rect 7477 8730 7483 8732
rect 7539 8730 7563 8732
rect 7619 8730 7643 8732
rect 7699 8730 7723 8732
rect 7779 8730 7785 8732
rect 7539 8678 7541 8730
rect 7721 8678 7723 8730
rect 7477 8676 7483 8678
rect 7539 8676 7563 8678
rect 7619 8676 7643 8678
rect 7699 8676 7723 8678
rect 7779 8676 7785 8678
rect 7477 8656 7785 8676
rect 9876 8498 9904 9318
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 10046 8392 10102 8401
rect 10046 8327 10048 8336
rect 10100 8327 10102 8336
rect 10048 8298 10100 8304
rect 9109 8188 9417 8208
rect 9109 8186 9115 8188
rect 9171 8186 9195 8188
rect 9251 8186 9275 8188
rect 9331 8186 9355 8188
rect 9411 8186 9417 8188
rect 9171 8134 9173 8186
rect 9353 8134 9355 8186
rect 9109 8132 9115 8134
rect 9171 8132 9195 8134
rect 9251 8132 9275 8134
rect 9331 8132 9355 8134
rect 9411 8132 9417 8134
rect 9109 8112 9417 8132
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 7477 7644 7785 7664
rect 7477 7642 7483 7644
rect 7539 7642 7563 7644
rect 7619 7642 7643 7644
rect 7699 7642 7723 7644
rect 7779 7642 7785 7644
rect 7539 7590 7541 7642
rect 7721 7590 7723 7642
rect 7477 7588 7483 7590
rect 7539 7588 7563 7590
rect 7619 7588 7643 7590
rect 7699 7588 7723 7590
rect 7779 7588 7785 7590
rect 7477 7568 7785 7588
rect 9876 7410 9904 7686
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 10046 7304 10102 7313
rect 10046 7239 10048 7248
rect 10100 7239 10102 7248
rect 10048 7210 10100 7216
rect 9109 7100 9417 7120
rect 9109 7098 9115 7100
rect 9171 7098 9195 7100
rect 9251 7098 9275 7100
rect 9331 7098 9355 7100
rect 9411 7098 9417 7100
rect 9171 7046 9173 7098
rect 9353 7046 9355 7098
rect 9109 7044 9115 7046
rect 9171 7044 9195 7046
rect 9251 7044 9275 7046
rect 9331 7044 9355 7046
rect 9411 7044 9417 7046
rect 9109 7024 9417 7044
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 7477 6556 7785 6576
rect 7477 6554 7483 6556
rect 7539 6554 7563 6556
rect 7619 6554 7643 6556
rect 7699 6554 7723 6556
rect 7779 6554 7785 6556
rect 7539 6502 7541 6554
rect 7721 6502 7723 6554
rect 7477 6500 7483 6502
rect 7539 6500 7563 6502
rect 7619 6500 7643 6502
rect 7699 6500 7723 6502
rect 7779 6500 7785 6502
rect 7477 6480 7785 6500
rect 9876 6322 9904 6598
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 6828 6180 6880 6186
rect 6828 6122 6880 6128
rect 9772 6112 9824 6118
rect 10048 6112 10100 6118
rect 9772 6054 9824 6060
rect 10046 6080 10048 6089
rect 10100 6080 10102 6089
rect 5845 6012 6153 6032
rect 5845 6010 5851 6012
rect 5907 6010 5931 6012
rect 5987 6010 6011 6012
rect 6067 6010 6091 6012
rect 6147 6010 6153 6012
rect 5907 5958 5909 6010
rect 6089 5958 6091 6010
rect 5845 5956 5851 5958
rect 5907 5956 5931 5958
rect 5987 5956 6011 5958
rect 6067 5956 6091 5958
rect 6147 5956 6153 5958
rect 5845 5936 6153 5956
rect 9109 6012 9417 6032
rect 9109 6010 9115 6012
rect 9171 6010 9195 6012
rect 9251 6010 9275 6012
rect 9331 6010 9355 6012
rect 9411 6010 9417 6012
rect 9171 5958 9173 6010
rect 9353 5958 9355 6010
rect 9109 5956 9115 5958
rect 9171 5956 9195 5958
rect 9251 5956 9275 5958
rect 9331 5956 9355 5958
rect 9411 5956 9417 5958
rect 9109 5936 9417 5956
rect 5080 5704 5132 5710
rect 5356 5704 5408 5710
rect 5132 5652 5356 5658
rect 5080 5646 5408 5652
rect 5092 5630 5396 5646
rect 4213 5468 4521 5488
rect 4213 5466 4219 5468
rect 4275 5466 4299 5468
rect 4355 5466 4379 5468
rect 4435 5466 4459 5468
rect 4515 5466 4521 5468
rect 4275 5414 4277 5466
rect 4457 5414 4459 5466
rect 4213 5412 4219 5414
rect 4275 5412 4299 5414
rect 4355 5412 4379 5414
rect 4435 5412 4459 5414
rect 4515 5412 4521 5414
rect 4213 5392 4521 5412
rect 5092 5234 5120 5630
rect 7477 5468 7785 5488
rect 7477 5466 7483 5468
rect 7539 5466 7563 5468
rect 7619 5466 7643 5468
rect 7699 5466 7723 5468
rect 7779 5466 7785 5468
rect 7539 5414 7541 5466
rect 7721 5414 7723 5466
rect 7477 5412 7483 5414
rect 7539 5412 7563 5414
rect 7619 5412 7643 5414
rect 7699 5412 7723 5414
rect 7779 5412 7785 5414
rect 7477 5392 7785 5412
rect 9784 5234 9812 6054
rect 10046 6015 10102 6024
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 4213 4380 4521 4400
rect 4213 4378 4219 4380
rect 4275 4378 4299 4380
rect 4355 4378 4379 4380
rect 4435 4378 4459 4380
rect 4515 4378 4521 4380
rect 4275 4326 4277 4378
rect 4457 4326 4459 4378
rect 4213 4324 4219 4326
rect 4275 4324 4299 4326
rect 4355 4324 4379 4326
rect 4435 4324 4459 4326
rect 4515 4324 4521 4326
rect 4213 4304 4521 4324
rect 4816 4214 4844 4966
rect 5845 4924 6153 4944
rect 5845 4922 5851 4924
rect 5907 4922 5931 4924
rect 5987 4922 6011 4924
rect 6067 4922 6091 4924
rect 6147 4922 6153 4924
rect 5907 4870 5909 4922
rect 6089 4870 6091 4922
rect 5845 4868 5851 4870
rect 5907 4868 5931 4870
rect 5987 4868 6011 4870
rect 6067 4868 6091 4870
rect 6147 4868 6153 4870
rect 5845 4848 6153 4868
rect 9109 4924 9417 4944
rect 9109 4922 9115 4924
rect 9171 4922 9195 4924
rect 9251 4922 9275 4924
rect 9331 4922 9355 4924
rect 9411 4922 9417 4924
rect 9171 4870 9173 4922
rect 9353 4870 9355 4922
rect 9109 4868 9115 4870
rect 9171 4868 9195 4870
rect 9251 4868 9275 4870
rect 9331 4868 9355 4870
rect 9411 4868 9417 4870
rect 9109 4848 9417 4868
rect 7477 4380 7785 4400
rect 7477 4378 7483 4380
rect 7539 4378 7563 4380
rect 7619 4378 7643 4380
rect 7699 4378 7723 4380
rect 7779 4378 7785 4380
rect 7539 4326 7541 4378
rect 7721 4326 7723 4378
rect 7477 4324 7483 4326
rect 7539 4324 7563 4326
rect 7619 4324 7643 4326
rect 7699 4324 7723 4326
rect 7779 4324 7785 4326
rect 7477 4304 7785 4324
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 5845 3836 6153 3856
rect 5845 3834 5851 3836
rect 5907 3834 5931 3836
rect 5987 3834 6011 3836
rect 6067 3834 6091 3836
rect 6147 3834 6153 3836
rect 5907 3782 5909 3834
rect 6089 3782 6091 3834
rect 5845 3780 5851 3782
rect 5907 3780 5931 3782
rect 5987 3780 6011 3782
rect 6067 3780 6091 3782
rect 6147 3780 6153 3782
rect 5845 3760 6153 3780
rect 9109 3836 9417 3856
rect 9109 3834 9115 3836
rect 9171 3834 9195 3836
rect 9251 3834 9275 3836
rect 9331 3834 9355 3836
rect 9411 3834 9417 3836
rect 9171 3782 9173 3834
rect 9353 3782 9355 3834
rect 9109 3780 9115 3782
rect 9171 3780 9195 3782
rect 9251 3780 9275 3782
rect 9331 3780 9355 3782
rect 9411 3780 9417 3782
rect 9109 3760 9417 3780
rect 9876 3534 9904 5510
rect 10048 5024 10100 5030
rect 10046 4992 10048 5001
rect 10100 4992 10102 5001
rect 10046 4927 10102 4936
rect 10048 3936 10100 3942
rect 10046 3904 10048 3913
rect 10100 3904 10102 3913
rect 10046 3839 10102 3848
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 4213 3292 4521 3312
rect 4213 3290 4219 3292
rect 4275 3290 4299 3292
rect 4355 3290 4379 3292
rect 4435 3290 4459 3292
rect 4515 3290 4521 3292
rect 4275 3238 4277 3290
rect 4457 3238 4459 3290
rect 4213 3236 4219 3238
rect 4275 3236 4299 3238
rect 4355 3236 4379 3238
rect 4435 3236 4459 3238
rect 4515 3236 4521 3238
rect 4213 3216 4521 3236
rect 7477 3292 7785 3312
rect 7477 3290 7483 3292
rect 7539 3290 7563 3292
rect 7619 3290 7643 3292
rect 7699 3290 7723 3292
rect 7779 3290 7785 3292
rect 7539 3238 7541 3290
rect 7721 3238 7723 3290
rect 7477 3236 7483 3238
rect 7539 3236 7563 3238
rect 7619 3236 7643 3238
rect 7699 3236 7723 3238
rect 7779 3236 7785 3238
rect 7477 3216 7785 3236
rect 10060 2825 10088 3334
rect 2582 2748 2890 2768
rect 2582 2746 2588 2748
rect 2644 2746 2668 2748
rect 2724 2746 2748 2748
rect 2804 2746 2828 2748
rect 2884 2746 2890 2748
rect 2644 2694 2646 2746
rect 2826 2694 2828 2746
rect 2582 2692 2588 2694
rect 2644 2692 2668 2694
rect 2724 2692 2748 2694
rect 2804 2692 2828 2694
rect 2884 2692 2890 2694
rect 2582 2672 2890 2692
rect 2976 2746 3096 2774
rect 10046 2816 10102 2825
rect 5845 2748 6153 2768
rect 5845 2746 5851 2748
rect 5907 2746 5931 2748
rect 5987 2746 6011 2748
rect 6067 2746 6091 2748
rect 6147 2746 6153 2748
rect 2976 2650 3004 2746
rect 5907 2694 5909 2746
rect 6089 2694 6091 2746
rect 5845 2692 5851 2694
rect 5907 2692 5931 2694
rect 5987 2692 6011 2694
rect 6067 2692 6091 2694
rect 6147 2692 6153 2694
rect 5845 2672 6153 2692
rect 9109 2748 9417 2768
rect 10046 2751 10102 2760
rect 9109 2746 9115 2748
rect 9171 2746 9195 2748
rect 9251 2746 9275 2748
rect 9331 2746 9355 2748
rect 9411 2746 9417 2748
rect 9171 2694 9173 2746
rect 9353 2694 9355 2746
rect 9109 2692 9115 2694
rect 9171 2692 9195 2694
rect 9251 2692 9275 2694
rect 9331 2692 9355 2694
rect 9411 2692 9417 2694
rect 9109 2672 9417 2692
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 2044 2440 2096 2446
rect 1308 2382 1360 2388
rect 1398 2408 1454 2417
rect 1320 1465 1348 2382
rect 2044 2382 2096 2388
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 1398 2343 1454 2352
rect 1306 1456 1362 1465
rect 1306 1391 1362 1400
rect 2056 1057 2084 2382
rect 2792 2009 2820 2382
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 4213 2204 4521 2224
rect 4213 2202 4219 2204
rect 4275 2202 4299 2204
rect 4355 2202 4379 2204
rect 4435 2202 4459 2204
rect 4515 2202 4521 2204
rect 4275 2150 4277 2202
rect 4457 2150 4459 2202
rect 4213 2148 4219 2150
rect 4275 2148 4299 2150
rect 4355 2148 4379 2150
rect 4435 2148 4459 2150
rect 4515 2148 4521 2150
rect 4213 2128 4521 2148
rect 7477 2204 7785 2224
rect 7477 2202 7483 2204
rect 7539 2202 7563 2204
rect 7619 2202 7643 2204
rect 7699 2202 7723 2204
rect 7779 2202 7785 2204
rect 7539 2150 7541 2202
rect 7721 2150 7723 2202
rect 7477 2148 7483 2150
rect 7539 2148 7563 2150
rect 7619 2148 7643 2150
rect 7699 2148 7723 2150
rect 7779 2148 7785 2150
rect 7477 2128 7785 2148
rect 2778 2000 2834 2009
rect 2778 1935 2834 1944
rect 10060 1737 10088 2246
rect 10046 1728 10102 1737
rect 10046 1663 10102 1672
rect 2042 1048 2098 1057
rect 2042 983 2098 992
rect 10968 672 11020 678
rect 10966 640 10968 649
rect 11020 640 11022 649
rect 10966 575 11022 584
<< via2 >>
rect 3146 79600 3202 79656
rect 3054 79192 3110 79248
rect 2962 78240 3018 78296
rect 2588 77818 2644 77820
rect 2668 77818 2724 77820
rect 2748 77818 2804 77820
rect 2828 77818 2884 77820
rect 2588 77766 2634 77818
rect 2634 77766 2644 77818
rect 2668 77766 2698 77818
rect 2698 77766 2710 77818
rect 2710 77766 2724 77818
rect 2748 77766 2762 77818
rect 2762 77766 2774 77818
rect 2774 77766 2804 77818
rect 2828 77766 2838 77818
rect 2838 77766 2884 77818
rect 2588 77764 2644 77766
rect 2668 77764 2724 77766
rect 2748 77764 2804 77766
rect 2828 77764 2884 77766
rect 2870 77560 2926 77616
rect 2042 77460 2044 77480
rect 2044 77460 2096 77480
rect 2096 77460 2098 77480
rect 2042 77424 2098 77460
rect 1490 76472 1546 76528
rect 1398 76064 1454 76120
rect 1306 75112 1362 75168
rect 1398 74296 1454 74352
rect 1306 73344 1362 73400
rect 1398 72936 1454 72992
rect 1306 71984 1362 72040
rect 1214 71576 1270 71632
rect 1398 71032 1454 71088
rect 1306 70216 1362 70272
rect 1214 69264 1270 69320
rect 1398 68856 1454 68912
rect 1306 68448 1362 68504
rect 2042 76880 2098 76936
rect 1674 70488 1730 70544
rect 1398 67904 1454 67960
rect 1490 67768 1546 67824
rect 1398 67496 1454 67552
rect 1398 66136 1454 66192
rect 1490 63416 1546 63472
rect 1398 62600 1454 62656
rect 1490 62056 1546 62112
rect 1398 61240 1454 61296
rect 1490 60696 1546 60752
rect 1398 60288 1454 60344
rect 1490 59880 1546 59936
rect 1398 58928 1454 58984
rect 2226 75520 2282 75576
rect 2042 72392 2098 72448
rect 1674 67088 1730 67144
rect 1490 58112 1546 58168
rect 1490 55800 1546 55856
rect 1490 55392 1546 55448
rect 1398 55256 1454 55312
rect 1490 54440 1546 54496
rect 1398 53624 1454 53680
rect 1490 52672 1546 52728
rect 1674 58248 1730 58304
rect 1398 51720 1454 51776
rect 1306 51176 1362 51232
rect 1950 65728 2006 65784
rect 1950 65184 2006 65240
rect 1950 62056 2006 62112
rect 2588 76730 2644 76732
rect 2668 76730 2724 76732
rect 2748 76730 2804 76732
rect 2828 76730 2884 76732
rect 2588 76678 2634 76730
rect 2634 76678 2644 76730
rect 2668 76678 2698 76730
rect 2698 76678 2710 76730
rect 2710 76678 2724 76730
rect 2748 76678 2762 76730
rect 2762 76678 2774 76730
rect 2774 76678 2804 76730
rect 2828 76678 2838 76730
rect 2838 76678 2884 76730
rect 2588 76676 2644 76678
rect 2668 76676 2724 76678
rect 2748 76676 2804 76678
rect 2828 76676 2884 76678
rect 2588 75642 2644 75644
rect 2668 75642 2724 75644
rect 2748 75642 2804 75644
rect 2828 75642 2884 75644
rect 2588 75590 2634 75642
rect 2634 75590 2644 75642
rect 2668 75590 2698 75642
rect 2698 75590 2710 75642
rect 2710 75590 2724 75642
rect 2748 75590 2762 75642
rect 2762 75590 2774 75642
rect 2774 75590 2804 75642
rect 2828 75590 2838 75642
rect 2838 75590 2884 75642
rect 2588 75588 2644 75590
rect 2668 75588 2724 75590
rect 2748 75588 2804 75590
rect 2828 75588 2884 75590
rect 9494 79328 9550 79384
rect 3974 78784 4030 78840
rect 5851 77818 5907 77820
rect 5931 77818 5987 77820
rect 6011 77818 6067 77820
rect 6091 77818 6147 77820
rect 5851 77766 5897 77818
rect 5897 77766 5907 77818
rect 5931 77766 5961 77818
rect 5961 77766 5973 77818
rect 5973 77766 5987 77818
rect 6011 77766 6025 77818
rect 6025 77766 6037 77818
rect 6037 77766 6067 77818
rect 6091 77766 6101 77818
rect 6101 77766 6147 77818
rect 5851 77764 5907 77766
rect 5931 77764 5987 77766
rect 6011 77764 6067 77766
rect 6091 77764 6147 77766
rect 9115 77818 9171 77820
rect 9195 77818 9251 77820
rect 9275 77818 9331 77820
rect 9355 77818 9411 77820
rect 9115 77766 9161 77818
rect 9161 77766 9171 77818
rect 9195 77766 9225 77818
rect 9225 77766 9237 77818
rect 9237 77766 9251 77818
rect 9275 77766 9289 77818
rect 9289 77766 9301 77818
rect 9301 77766 9331 77818
rect 9355 77766 9365 77818
rect 9365 77766 9411 77818
rect 9115 77764 9171 77766
rect 9195 77764 9251 77766
rect 9275 77764 9331 77766
rect 9355 77764 9411 77766
rect 10966 78260 11022 78296
rect 10966 78240 10968 78260
rect 10968 78240 11020 78260
rect 11020 78240 11022 78260
rect 4219 77274 4275 77276
rect 4299 77274 4355 77276
rect 4379 77274 4435 77276
rect 4459 77274 4515 77276
rect 4219 77222 4265 77274
rect 4265 77222 4275 77274
rect 4299 77222 4329 77274
rect 4329 77222 4341 77274
rect 4341 77222 4355 77274
rect 4379 77222 4393 77274
rect 4393 77222 4405 77274
rect 4405 77222 4435 77274
rect 4459 77222 4469 77274
rect 4469 77222 4515 77274
rect 4219 77220 4275 77222
rect 4299 77220 4355 77222
rect 4379 77220 4435 77222
rect 4459 77220 4515 77222
rect 2778 74704 2834 74760
rect 2588 74554 2644 74556
rect 2668 74554 2724 74556
rect 2748 74554 2804 74556
rect 2828 74554 2884 74556
rect 2588 74502 2634 74554
rect 2634 74502 2644 74554
rect 2668 74502 2698 74554
rect 2698 74502 2710 74554
rect 2710 74502 2724 74554
rect 2748 74502 2762 74554
rect 2762 74502 2774 74554
rect 2774 74502 2804 74554
rect 2828 74502 2838 74554
rect 2838 74502 2884 74554
rect 2588 74500 2644 74502
rect 2668 74500 2724 74502
rect 2748 74500 2804 74502
rect 2828 74500 2884 74502
rect 2870 73752 2926 73808
rect 2318 68992 2374 69048
rect 2226 68584 2282 68640
rect 2318 64812 2320 64832
rect 2320 64812 2372 64832
rect 2372 64812 2374 64832
rect 2318 64776 2374 64812
rect 2588 73466 2644 73468
rect 2668 73466 2724 73468
rect 2748 73466 2804 73468
rect 2828 73466 2884 73468
rect 2588 73414 2634 73466
rect 2634 73414 2644 73466
rect 2668 73414 2698 73466
rect 2698 73414 2710 73466
rect 2710 73414 2724 73466
rect 2748 73414 2762 73466
rect 2762 73414 2774 73466
rect 2774 73414 2804 73466
rect 2828 73414 2838 73466
rect 2838 73414 2884 73466
rect 2588 73412 2644 73414
rect 2668 73412 2724 73414
rect 2748 73412 2804 73414
rect 2828 73412 2884 73414
rect 2588 72378 2644 72380
rect 2668 72378 2724 72380
rect 2748 72378 2804 72380
rect 2828 72378 2884 72380
rect 2588 72326 2634 72378
rect 2634 72326 2644 72378
rect 2668 72326 2698 72378
rect 2698 72326 2710 72378
rect 2710 72326 2724 72378
rect 2748 72326 2762 72378
rect 2762 72326 2774 72378
rect 2774 72326 2804 72378
rect 2828 72326 2838 72378
rect 2838 72326 2884 72378
rect 2588 72324 2644 72326
rect 2668 72324 2724 72326
rect 2748 72324 2804 72326
rect 2828 72324 2884 72326
rect 2588 71290 2644 71292
rect 2668 71290 2724 71292
rect 2748 71290 2804 71292
rect 2828 71290 2884 71292
rect 2588 71238 2634 71290
rect 2634 71238 2644 71290
rect 2668 71238 2698 71290
rect 2698 71238 2710 71290
rect 2710 71238 2724 71290
rect 2748 71238 2762 71290
rect 2762 71238 2774 71290
rect 2774 71238 2804 71290
rect 2828 71238 2838 71290
rect 2838 71238 2884 71290
rect 2588 71236 2644 71238
rect 2668 71236 2724 71238
rect 2748 71236 2804 71238
rect 2828 71236 2884 71238
rect 2778 70624 2834 70680
rect 2588 70202 2644 70204
rect 2668 70202 2724 70204
rect 2748 70202 2804 70204
rect 2828 70202 2884 70204
rect 2588 70150 2634 70202
rect 2634 70150 2644 70202
rect 2668 70150 2698 70202
rect 2698 70150 2710 70202
rect 2710 70150 2724 70202
rect 2748 70150 2762 70202
rect 2762 70150 2774 70202
rect 2774 70150 2804 70202
rect 2828 70150 2838 70202
rect 2838 70150 2884 70202
rect 2588 70148 2644 70150
rect 2668 70148 2724 70150
rect 2748 70148 2804 70150
rect 2828 70148 2884 70150
rect 2870 69844 2872 69864
rect 2872 69844 2924 69864
rect 2924 69844 2926 69864
rect 2870 69808 2926 69844
rect 2588 69114 2644 69116
rect 2668 69114 2724 69116
rect 2748 69114 2804 69116
rect 2828 69114 2884 69116
rect 2588 69062 2634 69114
rect 2634 69062 2644 69114
rect 2668 69062 2698 69114
rect 2698 69062 2710 69114
rect 2710 69062 2724 69114
rect 2748 69062 2762 69114
rect 2762 69062 2774 69114
rect 2774 69062 2804 69114
rect 2828 69062 2838 69114
rect 2838 69062 2884 69114
rect 2588 69060 2644 69062
rect 2668 69060 2724 69062
rect 2748 69060 2804 69062
rect 2828 69060 2884 69062
rect 2588 68026 2644 68028
rect 2668 68026 2724 68028
rect 2748 68026 2804 68028
rect 2828 68026 2884 68028
rect 2588 67974 2634 68026
rect 2634 67974 2644 68026
rect 2668 67974 2698 68026
rect 2698 67974 2710 68026
rect 2710 67974 2724 68026
rect 2748 67974 2762 68026
rect 2762 67974 2774 68026
rect 2774 67974 2804 68026
rect 2828 67974 2838 68026
rect 2838 67974 2884 68026
rect 2588 67972 2644 67974
rect 2668 67972 2724 67974
rect 2748 67972 2804 67974
rect 2828 67972 2884 67974
rect 2588 66938 2644 66940
rect 2668 66938 2724 66940
rect 2748 66938 2804 66940
rect 2828 66938 2884 66940
rect 2588 66886 2634 66938
rect 2634 66886 2644 66938
rect 2668 66886 2698 66938
rect 2698 66886 2710 66938
rect 2710 66886 2724 66938
rect 2748 66886 2762 66938
rect 2762 66886 2774 66938
rect 2774 66886 2804 66938
rect 2828 66886 2838 66938
rect 2838 66886 2884 66938
rect 2588 66884 2644 66886
rect 2668 66884 2724 66886
rect 2748 66884 2804 66886
rect 2828 66884 2884 66886
rect 2778 66564 2834 66600
rect 2778 66544 2780 66564
rect 2780 66544 2832 66564
rect 2832 66544 2834 66564
rect 2588 65850 2644 65852
rect 2668 65850 2724 65852
rect 2748 65850 2804 65852
rect 2828 65850 2884 65852
rect 2588 65798 2634 65850
rect 2634 65798 2644 65850
rect 2668 65798 2698 65850
rect 2698 65798 2710 65850
rect 2710 65798 2724 65850
rect 2748 65798 2762 65850
rect 2762 65798 2774 65850
rect 2774 65798 2804 65850
rect 2828 65798 2838 65850
rect 2838 65798 2884 65850
rect 2588 65796 2644 65798
rect 2668 65796 2724 65798
rect 2748 65796 2804 65798
rect 2828 65796 2884 65798
rect 2588 64762 2644 64764
rect 2668 64762 2724 64764
rect 2748 64762 2804 64764
rect 2828 64762 2884 64764
rect 2588 64710 2634 64762
rect 2634 64710 2644 64762
rect 2668 64710 2698 64762
rect 2698 64710 2710 64762
rect 2710 64710 2724 64762
rect 2748 64710 2762 64762
rect 2762 64710 2774 64762
rect 2774 64710 2804 64762
rect 2828 64710 2838 64762
rect 2838 64710 2884 64762
rect 2588 64708 2644 64710
rect 2668 64708 2724 64710
rect 2748 64708 2804 64710
rect 2828 64708 2884 64710
rect 2588 63674 2644 63676
rect 2668 63674 2724 63676
rect 2748 63674 2804 63676
rect 2828 63674 2884 63676
rect 2588 63622 2634 63674
rect 2634 63622 2644 63674
rect 2668 63622 2698 63674
rect 2698 63622 2710 63674
rect 2710 63622 2724 63674
rect 2748 63622 2762 63674
rect 2762 63622 2774 63674
rect 2774 63622 2804 63674
rect 2828 63622 2838 63674
rect 2838 63622 2884 63674
rect 2588 63620 2644 63622
rect 2668 63620 2724 63622
rect 2748 63620 2804 63622
rect 2828 63620 2884 63622
rect 2226 61648 2282 61704
rect 2588 62586 2644 62588
rect 2668 62586 2724 62588
rect 2748 62586 2804 62588
rect 2828 62586 2884 62588
rect 2588 62534 2634 62586
rect 2634 62534 2644 62586
rect 2668 62534 2698 62586
rect 2698 62534 2710 62586
rect 2710 62534 2724 62586
rect 2748 62534 2762 62586
rect 2762 62534 2774 62586
rect 2774 62534 2804 62586
rect 2828 62534 2838 62586
rect 2838 62534 2884 62586
rect 2588 62532 2644 62534
rect 2668 62532 2724 62534
rect 2748 62532 2804 62534
rect 2828 62532 2884 62534
rect 2226 59492 2282 59528
rect 2226 59472 2228 59492
rect 2228 59472 2280 59492
rect 2280 59472 2282 59492
rect 2410 61512 2466 61568
rect 2042 53896 2098 53952
rect 1950 53352 2006 53408
rect 1582 51448 1638 51504
rect 1490 51312 1546 51368
rect 1582 51040 1638 51096
rect 1490 49136 1546 49192
rect 1490 48184 1546 48240
rect 1490 47776 1546 47832
rect 1950 51040 2006 51096
rect 1766 50224 1822 50280
rect 1490 46824 1546 46880
rect 1306 45464 1362 45520
rect 1490 46008 1546 46064
rect 1398 45056 1454 45112
rect 938 16768 994 16824
rect 1582 44784 1638 44840
rect 1490 44648 1546 44704
rect 1674 44240 1730 44296
rect 1582 44104 1638 44160
rect 1490 41928 1546 41984
rect 1398 41384 1454 41440
rect 1490 40976 1546 41032
rect 1490 40568 1546 40624
rect 1490 40160 1546 40216
rect 1490 39616 1546 39672
rect 1490 39244 1492 39264
rect 1492 39244 1544 39264
rect 1544 39244 1546 39264
rect 1490 39208 1546 39244
rect 1674 40296 1730 40352
rect 1490 38820 1546 38856
rect 1490 38800 1492 38820
rect 1492 38800 1544 38820
rect 1544 38800 1546 38820
rect 1398 38256 1454 38312
rect 1490 37848 1546 37904
rect 1858 44240 1914 44296
rect 1858 40024 1914 40080
rect 1582 36488 1638 36544
rect 1490 36080 1546 36136
rect 1582 35128 1638 35184
rect 1490 34720 1546 34776
rect 1582 34312 1638 34368
rect 1490 33768 1546 33824
rect 1582 33360 1638 33416
rect 1582 32988 1584 33008
rect 1584 32988 1636 33008
rect 1636 32988 1638 33008
rect 1582 32952 1638 32988
rect 1398 31048 1454 31104
rect 2318 56228 2374 56264
rect 2318 56208 2320 56228
rect 2320 56208 2372 56228
rect 2372 56208 2374 56228
rect 2226 55020 2228 55040
rect 2228 55020 2280 55040
rect 2280 55020 2282 55040
rect 2226 54984 2282 55020
rect 2226 54052 2282 54088
rect 2226 54032 2228 54052
rect 2228 54032 2280 54052
rect 2280 54032 2282 54052
rect 2226 53624 2282 53680
rect 2134 51312 2190 51368
rect 2318 53080 2374 53136
rect 2588 61498 2644 61500
rect 2668 61498 2724 61500
rect 2748 61498 2804 61500
rect 2828 61498 2884 61500
rect 2588 61446 2634 61498
rect 2634 61446 2644 61498
rect 2668 61446 2698 61498
rect 2698 61446 2710 61498
rect 2710 61446 2724 61498
rect 2748 61446 2762 61498
rect 2762 61446 2774 61498
rect 2774 61446 2804 61498
rect 2828 61446 2838 61498
rect 2838 61446 2884 61498
rect 2588 61444 2644 61446
rect 2668 61444 2724 61446
rect 2748 61444 2804 61446
rect 2828 61444 2884 61446
rect 2588 60410 2644 60412
rect 2668 60410 2724 60412
rect 2748 60410 2804 60412
rect 2828 60410 2884 60412
rect 2588 60358 2634 60410
rect 2634 60358 2644 60410
rect 2668 60358 2698 60410
rect 2698 60358 2710 60410
rect 2710 60358 2724 60410
rect 2748 60358 2762 60410
rect 2762 60358 2774 60410
rect 2774 60358 2804 60410
rect 2828 60358 2838 60410
rect 2838 60358 2884 60410
rect 2588 60356 2644 60358
rect 2668 60356 2724 60358
rect 2748 60356 2804 60358
rect 2828 60356 2884 60358
rect 2588 59322 2644 59324
rect 2668 59322 2724 59324
rect 2748 59322 2804 59324
rect 2828 59322 2884 59324
rect 2588 59270 2634 59322
rect 2634 59270 2644 59322
rect 2668 59270 2698 59322
rect 2698 59270 2710 59322
rect 2710 59270 2724 59322
rect 2748 59270 2762 59322
rect 2762 59270 2774 59322
rect 2774 59270 2804 59322
rect 2828 59270 2838 59322
rect 2838 59270 2884 59322
rect 2588 59268 2644 59270
rect 2668 59268 2724 59270
rect 2748 59268 2804 59270
rect 2828 59268 2884 59270
rect 2778 58520 2834 58576
rect 2588 58234 2644 58236
rect 2668 58234 2724 58236
rect 2748 58234 2804 58236
rect 2828 58234 2884 58236
rect 2588 58182 2634 58234
rect 2634 58182 2644 58234
rect 2668 58182 2698 58234
rect 2698 58182 2710 58234
rect 2710 58182 2724 58234
rect 2748 58182 2762 58234
rect 2762 58182 2774 58234
rect 2774 58182 2804 58234
rect 2828 58182 2838 58234
rect 2838 58182 2884 58234
rect 2588 58180 2644 58182
rect 2668 58180 2724 58182
rect 2748 58180 2804 58182
rect 2828 58180 2884 58182
rect 2502 57568 2558 57624
rect 2588 57146 2644 57148
rect 2668 57146 2724 57148
rect 2748 57146 2804 57148
rect 2828 57146 2884 57148
rect 2588 57094 2634 57146
rect 2634 57094 2644 57146
rect 2668 57094 2698 57146
rect 2698 57094 2710 57146
rect 2710 57094 2724 57146
rect 2748 57094 2762 57146
rect 2762 57094 2774 57146
rect 2774 57094 2804 57146
rect 2828 57094 2838 57146
rect 2838 57094 2884 57146
rect 2588 57092 2644 57094
rect 2668 57092 2724 57094
rect 2748 57092 2804 57094
rect 2828 57092 2884 57094
rect 2502 56752 2558 56808
rect 2588 56058 2644 56060
rect 2668 56058 2724 56060
rect 2748 56058 2804 56060
rect 2828 56058 2884 56060
rect 2588 56006 2634 56058
rect 2634 56006 2644 56058
rect 2668 56006 2698 56058
rect 2698 56006 2710 56058
rect 2710 56006 2724 56058
rect 2748 56006 2762 56058
rect 2762 56006 2774 56058
rect 2774 56006 2804 56058
rect 2828 56006 2838 56058
rect 2838 56006 2884 56058
rect 2588 56004 2644 56006
rect 2668 56004 2724 56006
rect 2748 56004 2804 56006
rect 2828 56004 2884 56006
rect 4219 76186 4275 76188
rect 4299 76186 4355 76188
rect 4379 76186 4435 76188
rect 4459 76186 4515 76188
rect 4219 76134 4265 76186
rect 4265 76134 4275 76186
rect 4299 76134 4329 76186
rect 4329 76134 4341 76186
rect 4341 76134 4355 76186
rect 4379 76134 4393 76186
rect 4393 76134 4405 76186
rect 4405 76134 4435 76186
rect 4459 76134 4469 76186
rect 4469 76134 4515 76186
rect 4219 76132 4275 76134
rect 4299 76132 4355 76134
rect 4379 76132 4435 76134
rect 4459 76132 4515 76134
rect 4219 75098 4275 75100
rect 4299 75098 4355 75100
rect 4379 75098 4435 75100
rect 4459 75098 4515 75100
rect 4219 75046 4265 75098
rect 4265 75046 4275 75098
rect 4299 75046 4329 75098
rect 4329 75046 4341 75098
rect 4341 75046 4355 75098
rect 4379 75046 4393 75098
rect 4393 75046 4405 75098
rect 4405 75046 4435 75098
rect 4459 75046 4469 75098
rect 4469 75046 4515 75098
rect 4219 75044 4275 75046
rect 4299 75044 4355 75046
rect 4379 75044 4435 75046
rect 4459 75044 4515 75046
rect 3146 64504 3202 64560
rect 3054 64368 3110 64424
rect 3146 57316 3202 57352
rect 3146 57296 3148 57316
rect 3148 57296 3200 57316
rect 3200 57296 3202 57316
rect 3054 56652 3056 56672
rect 3056 56652 3108 56672
rect 3108 56652 3110 56672
rect 3054 56616 3110 56652
rect 2588 54970 2644 54972
rect 2668 54970 2724 54972
rect 2748 54970 2804 54972
rect 2828 54970 2884 54972
rect 2588 54918 2634 54970
rect 2634 54918 2644 54970
rect 2668 54918 2698 54970
rect 2698 54918 2710 54970
rect 2710 54918 2724 54970
rect 2748 54918 2762 54970
rect 2762 54918 2774 54970
rect 2774 54918 2804 54970
rect 2828 54918 2838 54970
rect 2838 54918 2884 54970
rect 2588 54916 2644 54918
rect 2668 54916 2724 54918
rect 2748 54916 2804 54918
rect 2828 54916 2884 54918
rect 2588 53882 2644 53884
rect 2668 53882 2724 53884
rect 2748 53882 2804 53884
rect 2828 53882 2884 53884
rect 2588 53830 2634 53882
rect 2634 53830 2644 53882
rect 2668 53830 2698 53882
rect 2698 53830 2710 53882
rect 2710 53830 2724 53882
rect 2748 53830 2762 53882
rect 2762 53830 2774 53882
rect 2774 53830 2804 53882
rect 2828 53830 2838 53882
rect 2838 53830 2884 53882
rect 2588 53828 2644 53830
rect 2668 53828 2724 53830
rect 2748 53828 2804 53830
rect 2828 53828 2884 53830
rect 2318 51176 2374 51232
rect 2226 49580 2228 49600
rect 2228 49580 2280 49600
rect 2280 49580 2282 49600
rect 2226 49544 2282 49580
rect 2226 48612 2282 48648
rect 2226 48592 2228 48612
rect 2228 48592 2280 48612
rect 2280 48592 2282 48612
rect 2226 47232 2282 47288
rect 2226 45872 2282 45928
rect 2226 44784 2282 44840
rect 2226 42336 2282 42392
rect 2588 52794 2644 52796
rect 2668 52794 2724 52796
rect 2748 52794 2804 52796
rect 2828 52794 2884 52796
rect 2588 52742 2634 52794
rect 2634 52742 2644 52794
rect 2668 52742 2698 52794
rect 2698 52742 2710 52794
rect 2710 52742 2724 52794
rect 2748 52742 2762 52794
rect 2762 52742 2774 52794
rect 2774 52742 2804 52794
rect 2828 52742 2838 52794
rect 2838 52742 2884 52794
rect 2588 52740 2644 52742
rect 2668 52740 2724 52742
rect 2748 52740 2804 52742
rect 2828 52740 2884 52742
rect 2962 52264 3018 52320
rect 2588 51706 2644 51708
rect 2668 51706 2724 51708
rect 2748 51706 2804 51708
rect 2828 51706 2884 51708
rect 2588 51654 2634 51706
rect 2634 51654 2644 51706
rect 2668 51654 2698 51706
rect 2698 51654 2710 51706
rect 2710 51654 2724 51706
rect 2748 51654 2762 51706
rect 2762 51654 2774 51706
rect 2774 51654 2804 51706
rect 2828 51654 2838 51706
rect 2838 51654 2884 51706
rect 2588 51652 2644 51654
rect 2668 51652 2724 51654
rect 2748 51652 2804 51654
rect 2828 51652 2884 51654
rect 2962 50768 3018 50824
rect 2588 50618 2644 50620
rect 2668 50618 2724 50620
rect 2748 50618 2804 50620
rect 2828 50618 2884 50620
rect 2588 50566 2634 50618
rect 2634 50566 2644 50618
rect 2668 50566 2698 50618
rect 2698 50566 2710 50618
rect 2710 50566 2724 50618
rect 2748 50566 2762 50618
rect 2762 50566 2774 50618
rect 2774 50566 2804 50618
rect 2828 50566 2838 50618
rect 2838 50566 2884 50618
rect 2588 50564 2644 50566
rect 2668 50564 2724 50566
rect 2748 50564 2804 50566
rect 2828 50564 2884 50566
rect 2502 50224 2558 50280
rect 2502 49952 2558 50008
rect 3054 50632 3110 50688
rect 2588 49530 2644 49532
rect 2668 49530 2724 49532
rect 2748 49530 2804 49532
rect 2828 49530 2884 49532
rect 2588 49478 2634 49530
rect 2634 49478 2644 49530
rect 2668 49478 2698 49530
rect 2698 49478 2710 49530
rect 2710 49478 2724 49530
rect 2748 49478 2762 49530
rect 2762 49478 2774 49530
rect 2774 49478 2804 49530
rect 2828 49478 2838 49530
rect 2838 49478 2884 49530
rect 2588 49476 2644 49478
rect 2668 49476 2724 49478
rect 2748 49476 2804 49478
rect 2828 49476 2884 49478
rect 2588 48442 2644 48444
rect 2668 48442 2724 48444
rect 2748 48442 2804 48444
rect 2828 48442 2884 48444
rect 2588 48390 2634 48442
rect 2634 48390 2644 48442
rect 2668 48390 2698 48442
rect 2698 48390 2710 48442
rect 2710 48390 2724 48442
rect 2748 48390 2762 48442
rect 2762 48390 2774 48442
rect 2774 48390 2804 48442
rect 2828 48390 2838 48442
rect 2838 48390 2884 48442
rect 2588 48388 2644 48390
rect 2668 48388 2724 48390
rect 2748 48388 2804 48390
rect 2828 48388 2884 48390
rect 2870 47660 2926 47696
rect 2870 47640 2872 47660
rect 2872 47640 2924 47660
rect 2924 47640 2926 47660
rect 2588 47354 2644 47356
rect 2668 47354 2724 47356
rect 2748 47354 2804 47356
rect 2828 47354 2884 47356
rect 2588 47302 2634 47354
rect 2634 47302 2644 47354
rect 2668 47302 2698 47354
rect 2698 47302 2710 47354
rect 2710 47302 2724 47354
rect 2748 47302 2762 47354
rect 2762 47302 2774 47354
rect 2774 47302 2804 47354
rect 2828 47302 2838 47354
rect 2838 47302 2884 47354
rect 2588 47300 2644 47302
rect 2668 47300 2724 47302
rect 2748 47300 2804 47302
rect 2828 47300 2884 47302
rect 2502 46824 2558 46880
rect 2588 46266 2644 46268
rect 2668 46266 2724 46268
rect 2748 46266 2804 46268
rect 2828 46266 2884 46268
rect 2588 46214 2634 46266
rect 2634 46214 2644 46266
rect 2668 46214 2698 46266
rect 2698 46214 2710 46266
rect 2710 46214 2724 46266
rect 2748 46214 2762 46266
rect 2762 46214 2774 46266
rect 2774 46214 2804 46266
rect 2828 46214 2838 46266
rect 2838 46214 2884 46266
rect 2588 46212 2644 46214
rect 2668 46212 2724 46214
rect 2748 46212 2804 46214
rect 2828 46212 2884 46214
rect 2588 45178 2644 45180
rect 2668 45178 2724 45180
rect 2748 45178 2804 45180
rect 2828 45178 2884 45180
rect 2588 45126 2634 45178
rect 2634 45126 2644 45178
rect 2668 45126 2698 45178
rect 2698 45126 2710 45178
rect 2710 45126 2724 45178
rect 2748 45126 2762 45178
rect 2762 45126 2774 45178
rect 2774 45126 2804 45178
rect 2828 45126 2838 45178
rect 2838 45126 2884 45178
rect 2588 45124 2644 45126
rect 2668 45124 2724 45126
rect 2748 45124 2804 45126
rect 2828 45124 2884 45126
rect 3054 46436 3110 46472
rect 3054 46416 3056 46436
rect 3056 46416 3108 46436
rect 3108 46416 3110 46436
rect 2588 44090 2644 44092
rect 2668 44090 2724 44092
rect 2748 44090 2804 44092
rect 2828 44090 2884 44092
rect 2588 44038 2634 44090
rect 2634 44038 2644 44090
rect 2668 44038 2698 44090
rect 2698 44038 2710 44090
rect 2710 44038 2724 44090
rect 2748 44038 2762 44090
rect 2762 44038 2774 44090
rect 2774 44038 2804 44090
rect 2828 44038 2838 44090
rect 2838 44038 2884 44090
rect 2588 44036 2644 44038
rect 2668 44036 2724 44038
rect 2748 44036 2804 44038
rect 2828 44036 2884 44038
rect 2778 43288 2834 43344
rect 2588 43002 2644 43004
rect 2668 43002 2724 43004
rect 2748 43002 2804 43004
rect 2828 43002 2884 43004
rect 2588 42950 2634 43002
rect 2634 42950 2644 43002
rect 2668 42950 2698 43002
rect 2698 42950 2710 43002
rect 2710 42950 2724 43002
rect 2748 42950 2762 43002
rect 2762 42950 2774 43002
rect 2774 42950 2804 43002
rect 2828 42950 2838 43002
rect 2838 42950 2884 43002
rect 2588 42948 2644 42950
rect 2668 42948 2724 42950
rect 2748 42948 2804 42950
rect 2828 42948 2884 42950
rect 2502 42744 2558 42800
rect 2588 41914 2644 41916
rect 2668 41914 2724 41916
rect 2748 41914 2804 41916
rect 2828 41914 2884 41916
rect 2588 41862 2634 41914
rect 2634 41862 2644 41914
rect 2668 41862 2698 41914
rect 2698 41862 2710 41914
rect 2710 41862 2724 41914
rect 2748 41862 2762 41914
rect 2762 41862 2774 41914
rect 2774 41862 2804 41914
rect 2828 41862 2838 41914
rect 2838 41862 2884 41914
rect 2588 41860 2644 41862
rect 2668 41860 2724 41862
rect 2748 41860 2804 41862
rect 2828 41860 2884 41862
rect 2588 40826 2644 40828
rect 2668 40826 2724 40828
rect 2748 40826 2804 40828
rect 2828 40826 2884 40828
rect 2588 40774 2634 40826
rect 2634 40774 2644 40826
rect 2668 40774 2698 40826
rect 2698 40774 2710 40826
rect 2710 40774 2724 40826
rect 2748 40774 2762 40826
rect 2762 40774 2774 40826
rect 2774 40774 2804 40826
rect 2828 40774 2838 40826
rect 2838 40774 2884 40826
rect 2588 40772 2644 40774
rect 2668 40772 2724 40774
rect 2748 40772 2804 40774
rect 2828 40772 2884 40774
rect 2588 39738 2644 39740
rect 2668 39738 2724 39740
rect 2748 39738 2804 39740
rect 2828 39738 2884 39740
rect 2588 39686 2634 39738
rect 2634 39686 2644 39738
rect 2668 39686 2698 39738
rect 2698 39686 2710 39738
rect 2710 39686 2724 39738
rect 2748 39686 2762 39738
rect 2762 39686 2774 39738
rect 2774 39686 2804 39738
rect 2828 39686 2838 39738
rect 2838 39686 2884 39738
rect 2588 39684 2644 39686
rect 2668 39684 2724 39686
rect 2748 39684 2804 39686
rect 2828 39684 2884 39686
rect 2588 38650 2644 38652
rect 2668 38650 2724 38652
rect 2748 38650 2804 38652
rect 2828 38650 2884 38652
rect 2588 38598 2634 38650
rect 2634 38598 2644 38650
rect 2668 38598 2698 38650
rect 2698 38598 2710 38650
rect 2710 38598 2724 38650
rect 2748 38598 2762 38650
rect 2762 38598 2774 38650
rect 2774 38598 2804 38650
rect 2828 38598 2838 38650
rect 2838 38598 2884 38650
rect 2588 38596 2644 38598
rect 2668 38596 2724 38598
rect 2748 38596 2804 38598
rect 2828 38596 2884 38598
rect 2318 36896 2374 36952
rect 2318 36760 2374 36816
rect 2134 35808 2190 35864
rect 2588 37562 2644 37564
rect 2668 37562 2724 37564
rect 2748 37562 2804 37564
rect 2828 37562 2884 37564
rect 2588 37510 2634 37562
rect 2634 37510 2644 37562
rect 2668 37510 2698 37562
rect 2698 37510 2710 37562
rect 2710 37510 2724 37562
rect 2748 37510 2762 37562
rect 2762 37510 2774 37562
rect 2774 37510 2804 37562
rect 2828 37510 2838 37562
rect 2838 37510 2884 37562
rect 2588 37508 2644 37510
rect 2668 37508 2724 37510
rect 2748 37508 2804 37510
rect 2828 37508 2884 37510
rect 2588 36474 2644 36476
rect 2668 36474 2724 36476
rect 2748 36474 2804 36476
rect 2828 36474 2884 36476
rect 2588 36422 2634 36474
rect 2634 36422 2644 36474
rect 2668 36422 2698 36474
rect 2698 36422 2710 36474
rect 2710 36422 2724 36474
rect 2748 36422 2762 36474
rect 2762 36422 2774 36474
rect 2774 36422 2804 36474
rect 2828 36422 2838 36474
rect 2838 36422 2884 36474
rect 2588 36420 2644 36422
rect 2668 36420 2724 36422
rect 2748 36420 2804 36422
rect 2828 36420 2884 36422
rect 2594 35808 2650 35864
rect 2318 35556 2374 35592
rect 2318 35536 2320 35556
rect 2320 35536 2372 35556
rect 2372 35536 2374 35556
rect 2588 35386 2644 35388
rect 2668 35386 2724 35388
rect 2748 35386 2804 35388
rect 2828 35386 2884 35388
rect 2588 35334 2634 35386
rect 2634 35334 2644 35386
rect 2668 35334 2698 35386
rect 2698 35334 2710 35386
rect 2710 35334 2724 35386
rect 2748 35334 2762 35386
rect 2762 35334 2774 35386
rect 2774 35334 2804 35386
rect 2828 35334 2838 35386
rect 2838 35334 2884 35386
rect 2588 35332 2644 35334
rect 2668 35332 2724 35334
rect 2748 35332 2804 35334
rect 2828 35332 2884 35334
rect 2588 34298 2644 34300
rect 2668 34298 2724 34300
rect 2748 34298 2804 34300
rect 2828 34298 2884 34300
rect 2588 34246 2634 34298
rect 2634 34246 2644 34298
rect 2668 34246 2698 34298
rect 2698 34246 2710 34298
rect 2710 34246 2724 34298
rect 2748 34246 2762 34298
rect 2762 34246 2774 34298
rect 2774 34246 2804 34298
rect 2828 34246 2838 34298
rect 2838 34246 2884 34298
rect 2588 34244 2644 34246
rect 2668 34244 2724 34246
rect 2748 34244 2804 34246
rect 2828 34244 2884 34246
rect 2588 33210 2644 33212
rect 2668 33210 2724 33212
rect 2748 33210 2804 33212
rect 2828 33210 2884 33212
rect 2588 33158 2634 33210
rect 2634 33158 2644 33210
rect 2668 33158 2698 33210
rect 2698 33158 2710 33210
rect 2710 33158 2724 33210
rect 2748 33158 2762 33210
rect 2762 33158 2774 33210
rect 2774 33158 2804 33210
rect 2828 33158 2838 33210
rect 2838 33158 2884 33210
rect 2588 33156 2644 33158
rect 2668 33156 2724 33158
rect 2748 33156 2804 33158
rect 2828 33156 2884 33158
rect 2588 32122 2644 32124
rect 2668 32122 2724 32124
rect 2748 32122 2804 32124
rect 2828 32122 2884 32124
rect 2588 32070 2634 32122
rect 2634 32070 2644 32122
rect 2668 32070 2698 32122
rect 2698 32070 2710 32122
rect 2710 32070 2724 32122
rect 2748 32070 2762 32122
rect 2762 32070 2774 32122
rect 2774 32070 2804 32122
rect 2828 32070 2838 32122
rect 2838 32070 2884 32122
rect 2588 32068 2644 32070
rect 2668 32068 2724 32070
rect 2748 32068 2804 32070
rect 2828 32068 2884 32070
rect 2778 31592 2834 31648
rect 2588 31034 2644 31036
rect 2668 31034 2724 31036
rect 2748 31034 2804 31036
rect 2828 31034 2884 31036
rect 2588 30982 2634 31034
rect 2634 30982 2644 31034
rect 2668 30982 2698 31034
rect 2698 30982 2710 31034
rect 2710 30982 2724 31034
rect 2748 30982 2762 31034
rect 2762 30982 2774 31034
rect 2774 30982 2804 31034
rect 2828 30982 2838 31034
rect 2838 30982 2884 31034
rect 2588 30980 2644 30982
rect 2668 30980 2724 30982
rect 2748 30980 2804 30982
rect 2828 30980 2884 30982
rect 2778 30096 2834 30152
rect 2588 29946 2644 29948
rect 2668 29946 2724 29948
rect 2748 29946 2804 29948
rect 2828 29946 2884 29948
rect 2588 29894 2634 29946
rect 2634 29894 2644 29946
rect 2668 29894 2698 29946
rect 2698 29894 2710 29946
rect 2710 29894 2724 29946
rect 2748 29894 2762 29946
rect 2762 29894 2774 29946
rect 2774 29894 2804 29946
rect 2828 29894 2838 29946
rect 2838 29894 2884 29946
rect 2588 29892 2644 29894
rect 2668 29892 2724 29894
rect 2748 29892 2804 29894
rect 2828 29892 2884 29894
rect 2318 28872 2374 28928
rect 2588 28858 2644 28860
rect 2668 28858 2724 28860
rect 2748 28858 2804 28860
rect 2828 28858 2884 28860
rect 2588 28806 2634 28858
rect 2634 28806 2644 28858
rect 2668 28806 2698 28858
rect 2698 28806 2710 28858
rect 2710 28806 2724 28858
rect 2748 28806 2762 28858
rect 2762 28806 2774 28858
rect 2774 28806 2804 28858
rect 2828 28806 2838 28858
rect 2838 28806 2884 28858
rect 2588 28804 2644 28806
rect 2668 28804 2724 28806
rect 2748 28804 2804 28806
rect 2828 28804 2884 28806
rect 3606 55800 3662 55856
rect 3238 50768 3294 50824
rect 3422 50360 3478 50416
rect 3330 50224 3386 50280
rect 3238 49272 3294 49328
rect 3146 43152 3202 43208
rect 3238 37304 3294 37360
rect 4219 74010 4275 74012
rect 4299 74010 4355 74012
rect 4379 74010 4435 74012
rect 4459 74010 4515 74012
rect 4219 73958 4265 74010
rect 4265 73958 4275 74010
rect 4299 73958 4329 74010
rect 4329 73958 4341 74010
rect 4341 73958 4355 74010
rect 4379 73958 4393 74010
rect 4393 73958 4405 74010
rect 4405 73958 4435 74010
rect 4459 73958 4469 74010
rect 4469 73958 4515 74010
rect 4219 73956 4275 73958
rect 4299 73956 4355 73958
rect 4379 73956 4435 73958
rect 4459 73956 4515 73958
rect 4219 72922 4275 72924
rect 4299 72922 4355 72924
rect 4379 72922 4435 72924
rect 4459 72922 4515 72924
rect 4219 72870 4265 72922
rect 4265 72870 4275 72922
rect 4299 72870 4329 72922
rect 4329 72870 4341 72922
rect 4341 72870 4355 72922
rect 4379 72870 4393 72922
rect 4393 72870 4405 72922
rect 4405 72870 4435 72922
rect 4459 72870 4469 72922
rect 4469 72870 4515 72922
rect 4219 72868 4275 72870
rect 4299 72868 4355 72870
rect 4379 72868 4435 72870
rect 4459 72868 4515 72870
rect 4219 71834 4275 71836
rect 4299 71834 4355 71836
rect 4379 71834 4435 71836
rect 4459 71834 4515 71836
rect 4219 71782 4265 71834
rect 4265 71782 4275 71834
rect 4299 71782 4329 71834
rect 4329 71782 4341 71834
rect 4341 71782 4355 71834
rect 4379 71782 4393 71834
rect 4393 71782 4405 71834
rect 4405 71782 4435 71834
rect 4459 71782 4469 71834
rect 4469 71782 4515 71834
rect 4219 71780 4275 71782
rect 4299 71780 4355 71782
rect 4379 71780 4435 71782
rect 4459 71780 4515 71782
rect 4219 70746 4275 70748
rect 4299 70746 4355 70748
rect 4379 70746 4435 70748
rect 4459 70746 4515 70748
rect 4219 70694 4265 70746
rect 4265 70694 4275 70746
rect 4299 70694 4329 70746
rect 4329 70694 4341 70746
rect 4341 70694 4355 70746
rect 4379 70694 4393 70746
rect 4393 70694 4405 70746
rect 4405 70694 4435 70746
rect 4459 70694 4469 70746
rect 4469 70694 4515 70746
rect 4219 70692 4275 70694
rect 4299 70692 4355 70694
rect 4379 70692 4435 70694
rect 4459 70692 4515 70694
rect 4219 69658 4275 69660
rect 4299 69658 4355 69660
rect 4379 69658 4435 69660
rect 4459 69658 4515 69660
rect 4219 69606 4265 69658
rect 4265 69606 4275 69658
rect 4299 69606 4329 69658
rect 4329 69606 4341 69658
rect 4341 69606 4355 69658
rect 4379 69606 4393 69658
rect 4393 69606 4405 69658
rect 4405 69606 4435 69658
rect 4459 69606 4469 69658
rect 4469 69606 4515 69658
rect 4219 69604 4275 69606
rect 4299 69604 4355 69606
rect 4379 69604 4435 69606
rect 4459 69604 4515 69606
rect 4219 68570 4275 68572
rect 4299 68570 4355 68572
rect 4379 68570 4435 68572
rect 4459 68570 4515 68572
rect 4219 68518 4265 68570
rect 4265 68518 4275 68570
rect 4299 68518 4329 68570
rect 4329 68518 4341 68570
rect 4341 68518 4355 68570
rect 4379 68518 4393 68570
rect 4393 68518 4405 68570
rect 4405 68518 4435 68570
rect 4459 68518 4469 68570
rect 4469 68518 4515 68570
rect 4219 68516 4275 68518
rect 4299 68516 4355 68518
rect 4379 68516 4435 68518
rect 4459 68516 4515 68518
rect 7483 77274 7539 77276
rect 7563 77274 7619 77276
rect 7643 77274 7699 77276
rect 7723 77274 7779 77276
rect 7483 77222 7529 77274
rect 7529 77222 7539 77274
rect 7563 77222 7593 77274
rect 7593 77222 7605 77274
rect 7605 77222 7619 77274
rect 7643 77222 7657 77274
rect 7657 77222 7669 77274
rect 7669 77222 7699 77274
rect 7723 77222 7733 77274
rect 7733 77222 7779 77274
rect 7483 77220 7539 77222
rect 7563 77220 7619 77222
rect 7643 77220 7699 77222
rect 7723 77220 7779 77222
rect 5851 76730 5907 76732
rect 5931 76730 5987 76732
rect 6011 76730 6067 76732
rect 6091 76730 6147 76732
rect 5851 76678 5897 76730
rect 5897 76678 5907 76730
rect 5931 76678 5961 76730
rect 5961 76678 5973 76730
rect 5973 76678 5987 76730
rect 6011 76678 6025 76730
rect 6025 76678 6037 76730
rect 6037 76678 6067 76730
rect 6091 76678 6101 76730
rect 6101 76678 6147 76730
rect 5851 76676 5907 76678
rect 5931 76676 5987 76678
rect 6011 76676 6067 76678
rect 6091 76676 6147 76678
rect 9115 76730 9171 76732
rect 9195 76730 9251 76732
rect 9275 76730 9331 76732
rect 9355 76730 9411 76732
rect 9115 76678 9161 76730
rect 9161 76678 9171 76730
rect 9195 76678 9225 76730
rect 9225 76678 9237 76730
rect 9237 76678 9251 76730
rect 9275 76678 9289 76730
rect 9289 76678 9301 76730
rect 9301 76678 9331 76730
rect 9355 76678 9365 76730
rect 9365 76678 9411 76730
rect 9115 76676 9171 76678
rect 9195 76676 9251 76678
rect 9275 76676 9331 76678
rect 9355 76676 9411 76678
rect 7483 76186 7539 76188
rect 7563 76186 7619 76188
rect 7643 76186 7699 76188
rect 7723 76186 7779 76188
rect 7483 76134 7529 76186
rect 7529 76134 7539 76186
rect 7563 76134 7593 76186
rect 7593 76134 7605 76186
rect 7605 76134 7619 76186
rect 7643 76134 7657 76186
rect 7657 76134 7669 76186
rect 7669 76134 7699 76186
rect 7723 76134 7733 76186
rect 7733 76134 7779 76186
rect 7483 76132 7539 76134
rect 7563 76132 7619 76134
rect 7643 76132 7699 76134
rect 7723 76132 7779 76134
rect 5851 75642 5907 75644
rect 5931 75642 5987 75644
rect 6011 75642 6067 75644
rect 6091 75642 6147 75644
rect 5851 75590 5897 75642
rect 5897 75590 5907 75642
rect 5931 75590 5961 75642
rect 5961 75590 5973 75642
rect 5973 75590 5987 75642
rect 6011 75590 6025 75642
rect 6025 75590 6037 75642
rect 6037 75590 6067 75642
rect 6091 75590 6101 75642
rect 6101 75590 6147 75642
rect 5851 75588 5907 75590
rect 5931 75588 5987 75590
rect 6011 75588 6067 75590
rect 6091 75588 6147 75590
rect 9115 75642 9171 75644
rect 9195 75642 9251 75644
rect 9275 75642 9331 75644
rect 9355 75642 9411 75644
rect 9115 75590 9161 75642
rect 9161 75590 9171 75642
rect 9195 75590 9225 75642
rect 9225 75590 9237 75642
rect 9237 75590 9251 75642
rect 9275 75590 9289 75642
rect 9289 75590 9301 75642
rect 9301 75590 9331 75642
rect 9355 75590 9365 75642
rect 9365 75590 9411 75642
rect 9115 75588 9171 75590
rect 9195 75588 9251 75590
rect 9275 75588 9331 75590
rect 9355 75588 9411 75590
rect 7483 75098 7539 75100
rect 7563 75098 7619 75100
rect 7643 75098 7699 75100
rect 7723 75098 7779 75100
rect 7483 75046 7529 75098
rect 7529 75046 7539 75098
rect 7563 75046 7593 75098
rect 7593 75046 7605 75098
rect 7605 75046 7619 75098
rect 7643 75046 7657 75098
rect 7657 75046 7669 75098
rect 7669 75046 7699 75098
rect 7723 75046 7733 75098
rect 7733 75046 7779 75098
rect 7483 75044 7539 75046
rect 7563 75044 7619 75046
rect 7643 75044 7699 75046
rect 7723 75044 7779 75046
rect 10138 77152 10194 77208
rect 4219 67482 4275 67484
rect 4299 67482 4355 67484
rect 4379 67482 4435 67484
rect 4459 67482 4515 67484
rect 4219 67430 4265 67482
rect 4265 67430 4275 67482
rect 4299 67430 4329 67482
rect 4329 67430 4341 67482
rect 4341 67430 4355 67482
rect 4379 67430 4393 67482
rect 4393 67430 4405 67482
rect 4405 67430 4435 67482
rect 4459 67430 4469 67482
rect 4469 67430 4515 67482
rect 4219 67428 4275 67430
rect 4299 67428 4355 67430
rect 4379 67428 4435 67430
rect 4459 67428 4515 67430
rect 4219 66394 4275 66396
rect 4299 66394 4355 66396
rect 4379 66394 4435 66396
rect 4459 66394 4515 66396
rect 4219 66342 4265 66394
rect 4265 66342 4275 66394
rect 4299 66342 4329 66394
rect 4329 66342 4341 66394
rect 4341 66342 4355 66394
rect 4379 66342 4393 66394
rect 4393 66342 4405 66394
rect 4405 66342 4435 66394
rect 4459 66342 4469 66394
rect 4469 66342 4515 66394
rect 4219 66340 4275 66342
rect 4299 66340 4355 66342
rect 4379 66340 4435 66342
rect 4459 66340 4515 66342
rect 3974 63960 4030 64016
rect 3974 63008 4030 63064
rect 3974 54712 4030 54768
rect 3606 50768 3662 50824
rect 3790 51448 3846 51504
rect 4219 65306 4275 65308
rect 4299 65306 4355 65308
rect 4379 65306 4435 65308
rect 4459 65306 4515 65308
rect 4219 65254 4265 65306
rect 4265 65254 4275 65306
rect 4299 65254 4329 65306
rect 4329 65254 4341 65306
rect 4341 65254 4355 65306
rect 4379 65254 4393 65306
rect 4393 65254 4405 65306
rect 4405 65254 4435 65306
rect 4459 65254 4469 65306
rect 4469 65254 4515 65306
rect 4219 65252 4275 65254
rect 4299 65252 4355 65254
rect 4379 65252 4435 65254
rect 4459 65252 4515 65254
rect 4219 64218 4275 64220
rect 4299 64218 4355 64220
rect 4379 64218 4435 64220
rect 4459 64218 4515 64220
rect 4219 64166 4265 64218
rect 4265 64166 4275 64218
rect 4299 64166 4329 64218
rect 4329 64166 4341 64218
rect 4341 64166 4355 64218
rect 4379 64166 4393 64218
rect 4393 64166 4405 64218
rect 4405 64166 4435 64218
rect 4459 64166 4469 64218
rect 4469 64166 4515 64218
rect 4219 64164 4275 64166
rect 4299 64164 4355 64166
rect 4379 64164 4435 64166
rect 4459 64164 4515 64166
rect 4219 63130 4275 63132
rect 4299 63130 4355 63132
rect 4379 63130 4435 63132
rect 4459 63130 4515 63132
rect 4219 63078 4265 63130
rect 4265 63078 4275 63130
rect 4299 63078 4329 63130
rect 4329 63078 4341 63130
rect 4341 63078 4355 63130
rect 4379 63078 4393 63130
rect 4393 63078 4405 63130
rect 4405 63078 4435 63130
rect 4459 63078 4469 63130
rect 4469 63078 4515 63130
rect 4219 63076 4275 63078
rect 4299 63076 4355 63078
rect 4379 63076 4435 63078
rect 4459 63076 4515 63078
rect 4219 62042 4275 62044
rect 4299 62042 4355 62044
rect 4379 62042 4435 62044
rect 4459 62042 4515 62044
rect 4219 61990 4265 62042
rect 4265 61990 4275 62042
rect 4299 61990 4329 62042
rect 4329 61990 4341 62042
rect 4341 61990 4355 62042
rect 4379 61990 4393 62042
rect 4393 61990 4405 62042
rect 4405 61990 4435 62042
rect 4459 61990 4469 62042
rect 4469 61990 4515 62042
rect 4219 61988 4275 61990
rect 4299 61988 4355 61990
rect 4379 61988 4435 61990
rect 4459 61988 4515 61990
rect 4219 60954 4275 60956
rect 4299 60954 4355 60956
rect 4379 60954 4435 60956
rect 4459 60954 4515 60956
rect 4219 60902 4265 60954
rect 4265 60902 4275 60954
rect 4299 60902 4329 60954
rect 4329 60902 4341 60954
rect 4341 60902 4355 60954
rect 4379 60902 4393 60954
rect 4393 60902 4405 60954
rect 4405 60902 4435 60954
rect 4459 60902 4469 60954
rect 4469 60902 4515 60954
rect 4219 60900 4275 60902
rect 4299 60900 4355 60902
rect 4379 60900 4435 60902
rect 4459 60900 4515 60902
rect 4219 59866 4275 59868
rect 4299 59866 4355 59868
rect 4379 59866 4435 59868
rect 4459 59866 4515 59868
rect 4219 59814 4265 59866
rect 4265 59814 4275 59866
rect 4299 59814 4329 59866
rect 4329 59814 4341 59866
rect 4341 59814 4355 59866
rect 4379 59814 4393 59866
rect 4393 59814 4405 59866
rect 4405 59814 4435 59866
rect 4459 59814 4469 59866
rect 4469 59814 4515 59866
rect 4219 59812 4275 59814
rect 4299 59812 4355 59814
rect 4379 59812 4435 59814
rect 4459 59812 4515 59814
rect 4219 58778 4275 58780
rect 4299 58778 4355 58780
rect 4379 58778 4435 58780
rect 4459 58778 4515 58780
rect 4219 58726 4265 58778
rect 4265 58726 4275 58778
rect 4299 58726 4329 58778
rect 4329 58726 4341 58778
rect 4341 58726 4355 58778
rect 4379 58726 4393 58778
rect 4393 58726 4405 58778
rect 4405 58726 4435 58778
rect 4459 58726 4469 58778
rect 4469 58726 4515 58778
rect 4219 58724 4275 58726
rect 4299 58724 4355 58726
rect 4379 58724 4435 58726
rect 4459 58724 4515 58726
rect 4219 57690 4275 57692
rect 4299 57690 4355 57692
rect 4379 57690 4435 57692
rect 4459 57690 4515 57692
rect 4219 57638 4265 57690
rect 4265 57638 4275 57690
rect 4299 57638 4329 57690
rect 4329 57638 4341 57690
rect 4341 57638 4355 57690
rect 4379 57638 4393 57690
rect 4393 57638 4405 57690
rect 4405 57638 4435 57690
rect 4459 57638 4469 57690
rect 4469 57638 4515 57690
rect 4219 57636 4275 57638
rect 4299 57636 4355 57638
rect 4379 57636 4435 57638
rect 4459 57636 4515 57638
rect 4219 56602 4275 56604
rect 4299 56602 4355 56604
rect 4379 56602 4435 56604
rect 4459 56602 4515 56604
rect 4219 56550 4265 56602
rect 4265 56550 4275 56602
rect 4299 56550 4329 56602
rect 4329 56550 4341 56602
rect 4341 56550 4355 56602
rect 4379 56550 4393 56602
rect 4393 56550 4405 56602
rect 4405 56550 4435 56602
rect 4459 56550 4469 56602
rect 4469 56550 4515 56602
rect 4219 56548 4275 56550
rect 4299 56548 4355 56550
rect 4379 56548 4435 56550
rect 4459 56548 4515 56550
rect 4219 55514 4275 55516
rect 4299 55514 4355 55516
rect 4379 55514 4435 55516
rect 4459 55514 4515 55516
rect 4219 55462 4265 55514
rect 4265 55462 4275 55514
rect 4299 55462 4329 55514
rect 4329 55462 4341 55514
rect 4341 55462 4355 55514
rect 4379 55462 4393 55514
rect 4393 55462 4405 55514
rect 4405 55462 4435 55514
rect 4459 55462 4469 55514
rect 4469 55462 4515 55514
rect 4219 55460 4275 55462
rect 4299 55460 4355 55462
rect 4379 55460 4435 55462
rect 4459 55460 4515 55462
rect 4219 54426 4275 54428
rect 4299 54426 4355 54428
rect 4379 54426 4435 54428
rect 4459 54426 4515 54428
rect 4219 54374 4265 54426
rect 4265 54374 4275 54426
rect 4299 54374 4329 54426
rect 4329 54374 4341 54426
rect 4341 54374 4355 54426
rect 4379 54374 4393 54426
rect 4393 54374 4405 54426
rect 4405 54374 4435 54426
rect 4459 54374 4469 54426
rect 4469 54374 4515 54426
rect 4219 54372 4275 54374
rect 4299 54372 4355 54374
rect 4379 54372 4435 54374
rect 4459 54372 4515 54374
rect 4219 53338 4275 53340
rect 4299 53338 4355 53340
rect 4379 53338 4435 53340
rect 4459 53338 4515 53340
rect 4219 53286 4265 53338
rect 4265 53286 4275 53338
rect 4299 53286 4329 53338
rect 4329 53286 4341 53338
rect 4341 53286 4355 53338
rect 4379 53286 4393 53338
rect 4393 53286 4405 53338
rect 4405 53286 4435 53338
rect 4459 53286 4469 53338
rect 4469 53286 4515 53338
rect 4219 53284 4275 53286
rect 4299 53284 4355 53286
rect 4379 53284 4435 53286
rect 4459 53284 4515 53286
rect 3974 51032 4030 51088
rect 4802 56208 4858 56264
rect 4219 52250 4275 52252
rect 4299 52250 4355 52252
rect 4379 52250 4435 52252
rect 4459 52250 4515 52252
rect 4219 52198 4265 52250
rect 4265 52198 4275 52250
rect 4299 52198 4329 52250
rect 4329 52198 4341 52250
rect 4341 52198 4355 52250
rect 4379 52198 4393 52250
rect 4393 52198 4405 52250
rect 4405 52198 4435 52250
rect 4459 52198 4469 52250
rect 4469 52198 4515 52250
rect 4219 52196 4275 52198
rect 4299 52196 4355 52198
rect 4379 52196 4435 52198
rect 4459 52196 4515 52198
rect 4219 51162 4275 51164
rect 4299 51162 4355 51164
rect 4379 51162 4435 51164
rect 4459 51162 4515 51164
rect 4219 51110 4265 51162
rect 4265 51110 4275 51162
rect 4299 51110 4329 51162
rect 4329 51110 4341 51162
rect 4341 51110 4355 51162
rect 4379 51110 4393 51162
rect 4393 51110 4405 51162
rect 4405 51110 4435 51162
rect 4459 51110 4469 51162
rect 4469 51110 4515 51162
rect 4219 51108 4275 51110
rect 4299 51108 4355 51110
rect 4379 51108 4435 51110
rect 4459 51108 4515 51110
rect 3882 47640 3938 47696
rect 4219 50074 4275 50076
rect 4299 50074 4355 50076
rect 4379 50074 4435 50076
rect 4459 50074 4515 50076
rect 4219 50022 4265 50074
rect 4265 50022 4275 50074
rect 4299 50022 4329 50074
rect 4329 50022 4341 50074
rect 4341 50022 4355 50074
rect 4379 50022 4393 50074
rect 4393 50022 4405 50074
rect 4405 50022 4435 50074
rect 4459 50022 4469 50074
rect 4469 50022 4515 50074
rect 4219 50020 4275 50022
rect 4299 50020 4355 50022
rect 4379 50020 4435 50022
rect 4459 50020 4515 50022
rect 4219 48986 4275 48988
rect 4299 48986 4355 48988
rect 4379 48986 4435 48988
rect 4459 48986 4515 48988
rect 4219 48934 4265 48986
rect 4265 48934 4275 48986
rect 4299 48934 4329 48986
rect 4329 48934 4341 48986
rect 4341 48934 4355 48986
rect 4379 48934 4393 48986
rect 4393 48934 4405 48986
rect 4405 48934 4435 48986
rect 4459 48934 4469 48986
rect 4469 48934 4515 48986
rect 4219 48932 4275 48934
rect 4299 48932 4355 48934
rect 4379 48932 4435 48934
rect 4459 48932 4515 48934
rect 4434 48728 4490 48784
rect 4434 48184 4490 48240
rect 4526 48048 4582 48104
rect 4219 47898 4275 47900
rect 4299 47898 4355 47900
rect 4379 47898 4435 47900
rect 4459 47898 4515 47900
rect 4219 47846 4265 47898
rect 4265 47846 4275 47898
rect 4299 47846 4329 47898
rect 4329 47846 4341 47898
rect 4341 47846 4355 47898
rect 4379 47846 4393 47898
rect 4393 47846 4405 47898
rect 4405 47846 4435 47898
rect 4459 47846 4469 47898
rect 4469 47846 4515 47898
rect 4219 47844 4275 47846
rect 4299 47844 4355 47846
rect 4379 47844 4435 47846
rect 4459 47844 4515 47846
rect 4219 46810 4275 46812
rect 4299 46810 4355 46812
rect 4379 46810 4435 46812
rect 4459 46810 4515 46812
rect 4219 46758 4265 46810
rect 4265 46758 4275 46810
rect 4299 46758 4329 46810
rect 4329 46758 4341 46810
rect 4341 46758 4355 46810
rect 4379 46758 4393 46810
rect 4393 46758 4405 46810
rect 4405 46758 4435 46810
rect 4459 46758 4469 46810
rect 4469 46758 4515 46810
rect 4219 46756 4275 46758
rect 4299 46756 4355 46758
rect 4379 46756 4435 46758
rect 4459 46756 4515 46758
rect 4219 45722 4275 45724
rect 4299 45722 4355 45724
rect 4379 45722 4435 45724
rect 4459 45722 4515 45724
rect 4219 45670 4265 45722
rect 4265 45670 4275 45722
rect 4299 45670 4329 45722
rect 4329 45670 4341 45722
rect 4341 45670 4355 45722
rect 4379 45670 4393 45722
rect 4393 45670 4405 45722
rect 4405 45670 4435 45722
rect 4459 45670 4469 45722
rect 4469 45670 4515 45722
rect 4219 45668 4275 45670
rect 4299 45668 4355 45670
rect 4379 45668 4435 45670
rect 4459 45668 4515 45670
rect 4219 44634 4275 44636
rect 4299 44634 4355 44636
rect 4379 44634 4435 44636
rect 4459 44634 4515 44636
rect 4219 44582 4265 44634
rect 4265 44582 4275 44634
rect 4299 44582 4329 44634
rect 4329 44582 4341 44634
rect 4341 44582 4355 44634
rect 4379 44582 4393 44634
rect 4393 44582 4405 44634
rect 4405 44582 4435 44634
rect 4459 44582 4469 44634
rect 4469 44582 4515 44634
rect 4219 44580 4275 44582
rect 4299 44580 4355 44582
rect 4379 44580 4435 44582
rect 4459 44580 4515 44582
rect 3974 43696 4030 43752
rect 4219 43546 4275 43548
rect 4299 43546 4355 43548
rect 4379 43546 4435 43548
rect 4459 43546 4515 43548
rect 4219 43494 4265 43546
rect 4265 43494 4275 43546
rect 4299 43494 4329 43546
rect 4329 43494 4341 43546
rect 4341 43494 4355 43546
rect 4379 43494 4393 43546
rect 4393 43494 4405 43546
rect 4405 43494 4435 43546
rect 4459 43494 4469 43546
rect 4469 43494 4515 43546
rect 4219 43492 4275 43494
rect 4299 43492 4355 43494
rect 4379 43492 4435 43494
rect 4459 43492 4515 43494
rect 4219 42458 4275 42460
rect 4299 42458 4355 42460
rect 4379 42458 4435 42460
rect 4459 42458 4515 42460
rect 4219 42406 4265 42458
rect 4265 42406 4275 42458
rect 4299 42406 4329 42458
rect 4329 42406 4341 42458
rect 4341 42406 4355 42458
rect 4379 42406 4393 42458
rect 4393 42406 4405 42458
rect 4405 42406 4435 42458
rect 4459 42406 4469 42458
rect 4469 42406 4515 42458
rect 4219 42404 4275 42406
rect 4299 42404 4355 42406
rect 4379 42404 4435 42406
rect 4459 42404 4515 42406
rect 3054 32408 3110 32464
rect 3238 32272 3294 32328
rect 3146 30232 3202 30288
rect 3238 29280 3294 29336
rect 2588 27770 2644 27772
rect 2668 27770 2724 27772
rect 2748 27770 2804 27772
rect 2828 27770 2884 27772
rect 2588 27718 2634 27770
rect 2634 27718 2644 27770
rect 2668 27718 2698 27770
rect 2698 27718 2710 27770
rect 2710 27718 2724 27770
rect 2748 27718 2762 27770
rect 2762 27718 2774 27770
rect 2774 27718 2804 27770
rect 2828 27718 2838 27770
rect 2838 27718 2884 27770
rect 2588 27716 2644 27718
rect 2668 27716 2724 27718
rect 2748 27716 2804 27718
rect 2828 27716 2884 27718
rect 3054 27920 3110 27976
rect 3146 27512 3202 27568
rect 2226 27104 2282 27160
rect 2870 26832 2926 26888
rect 2588 26682 2644 26684
rect 2668 26682 2724 26684
rect 2748 26682 2804 26684
rect 2828 26682 2884 26684
rect 2588 26630 2634 26682
rect 2634 26630 2644 26682
rect 2668 26630 2698 26682
rect 2698 26630 2710 26682
rect 2710 26630 2724 26682
rect 2748 26630 2762 26682
rect 2762 26630 2774 26682
rect 2774 26630 2804 26682
rect 2828 26630 2838 26682
rect 2838 26630 2884 26682
rect 2588 26628 2644 26630
rect 2668 26628 2724 26630
rect 2748 26628 2804 26630
rect 2828 26628 2884 26630
rect 1398 24656 1454 24712
rect 1490 23432 1546 23488
rect 1490 23024 1546 23080
rect 2042 26152 2098 26208
rect 2226 25744 2282 25800
rect 2588 25594 2644 25596
rect 2668 25594 2724 25596
rect 2748 25594 2804 25596
rect 2828 25594 2884 25596
rect 2588 25542 2634 25594
rect 2634 25542 2644 25594
rect 2668 25542 2698 25594
rect 2698 25542 2710 25594
rect 2710 25542 2724 25594
rect 2748 25542 2762 25594
rect 2762 25542 2774 25594
rect 2774 25542 2804 25594
rect 2828 25542 2838 25594
rect 2838 25542 2884 25594
rect 2588 25540 2644 25542
rect 2668 25540 2724 25542
rect 2748 25540 2804 25542
rect 2828 25540 2884 25542
rect 2870 25236 2872 25256
rect 2872 25236 2924 25256
rect 2924 25236 2926 25256
rect 2870 25200 2926 25236
rect 2226 24792 2282 24848
rect 2588 24506 2644 24508
rect 2668 24506 2724 24508
rect 2748 24506 2804 24508
rect 2828 24506 2884 24508
rect 2588 24454 2634 24506
rect 2634 24454 2644 24506
rect 2668 24454 2698 24506
rect 2698 24454 2710 24506
rect 2710 24454 2724 24506
rect 2748 24454 2762 24506
rect 2762 24454 2774 24506
rect 2774 24454 2804 24506
rect 2828 24454 2838 24506
rect 2838 24454 2884 24506
rect 2588 24452 2644 24454
rect 2668 24452 2724 24454
rect 2748 24452 2804 24454
rect 2828 24452 2884 24454
rect 2870 23976 2926 24032
rect 2042 23568 2098 23624
rect 2588 23418 2644 23420
rect 2668 23418 2724 23420
rect 2748 23418 2804 23420
rect 2828 23418 2884 23420
rect 2588 23366 2634 23418
rect 2634 23366 2644 23418
rect 2668 23366 2698 23418
rect 2698 23366 2710 23418
rect 2710 23366 2724 23418
rect 2748 23366 2762 23418
rect 2762 23366 2774 23418
rect 2774 23366 2804 23418
rect 2828 23366 2838 23418
rect 2838 23366 2884 23418
rect 2588 23364 2644 23366
rect 2668 23364 2724 23366
rect 2748 23364 2804 23366
rect 2828 23364 2884 23366
rect 4219 41370 4275 41372
rect 4299 41370 4355 41372
rect 4379 41370 4435 41372
rect 4459 41370 4515 41372
rect 4219 41318 4265 41370
rect 4265 41318 4275 41370
rect 4299 41318 4329 41370
rect 4329 41318 4341 41370
rect 4341 41318 4355 41370
rect 4379 41318 4393 41370
rect 4393 41318 4405 41370
rect 4405 41318 4435 41370
rect 4459 41318 4469 41370
rect 4469 41318 4515 41370
rect 4219 41316 4275 41318
rect 4299 41316 4355 41318
rect 4379 41316 4435 41318
rect 4459 41316 4515 41318
rect 4219 40282 4275 40284
rect 4299 40282 4355 40284
rect 4379 40282 4435 40284
rect 4459 40282 4515 40284
rect 4219 40230 4265 40282
rect 4265 40230 4275 40282
rect 4299 40230 4329 40282
rect 4329 40230 4341 40282
rect 4341 40230 4355 40282
rect 4379 40230 4393 40282
rect 4393 40230 4405 40282
rect 4405 40230 4435 40282
rect 4459 40230 4469 40282
rect 4469 40230 4515 40282
rect 4219 40228 4275 40230
rect 4299 40228 4355 40230
rect 4379 40228 4435 40230
rect 4459 40228 4515 40230
rect 4219 39194 4275 39196
rect 4299 39194 4355 39196
rect 4379 39194 4435 39196
rect 4459 39194 4515 39196
rect 4219 39142 4265 39194
rect 4265 39142 4275 39194
rect 4299 39142 4329 39194
rect 4329 39142 4341 39194
rect 4341 39142 4355 39194
rect 4379 39142 4393 39194
rect 4393 39142 4405 39194
rect 4405 39142 4435 39194
rect 4459 39142 4469 39194
rect 4469 39142 4515 39194
rect 4219 39140 4275 39142
rect 4299 39140 4355 39142
rect 4379 39140 4435 39142
rect 4459 39140 4515 39142
rect 4219 38106 4275 38108
rect 4299 38106 4355 38108
rect 4379 38106 4435 38108
rect 4459 38106 4515 38108
rect 4219 38054 4265 38106
rect 4265 38054 4275 38106
rect 4299 38054 4329 38106
rect 4329 38054 4341 38106
rect 4341 38054 4355 38106
rect 4379 38054 4393 38106
rect 4393 38054 4405 38106
rect 4405 38054 4435 38106
rect 4459 38054 4469 38106
rect 4469 38054 4515 38106
rect 4219 38052 4275 38054
rect 4299 38052 4355 38054
rect 4379 38052 4435 38054
rect 4459 38052 4515 38054
rect 4219 37018 4275 37020
rect 4299 37018 4355 37020
rect 4379 37018 4435 37020
rect 4459 37018 4515 37020
rect 4219 36966 4265 37018
rect 4265 36966 4275 37018
rect 4299 36966 4329 37018
rect 4329 36966 4341 37018
rect 4341 36966 4355 37018
rect 4379 36966 4393 37018
rect 4393 36966 4405 37018
rect 4405 36966 4435 37018
rect 4459 36966 4469 37018
rect 4469 36966 4515 37018
rect 4219 36964 4275 36966
rect 4299 36964 4355 36966
rect 4379 36964 4435 36966
rect 4459 36964 4515 36966
rect 4219 35930 4275 35932
rect 4299 35930 4355 35932
rect 4379 35930 4435 35932
rect 4459 35930 4515 35932
rect 3974 30676 3976 30696
rect 3976 30676 4028 30696
rect 4028 30676 4030 30696
rect 3974 30640 4030 30676
rect 3514 28464 3570 28520
rect 4219 35878 4265 35930
rect 4265 35878 4275 35930
rect 4299 35878 4329 35930
rect 4329 35878 4341 35930
rect 4341 35878 4355 35930
rect 4379 35878 4393 35930
rect 4393 35878 4405 35930
rect 4405 35878 4435 35930
rect 4459 35878 4469 35930
rect 4469 35878 4515 35930
rect 4219 35876 4275 35878
rect 4299 35876 4355 35878
rect 4379 35876 4435 35878
rect 4459 35876 4515 35878
rect 4219 34842 4275 34844
rect 4299 34842 4355 34844
rect 4379 34842 4435 34844
rect 4459 34842 4515 34844
rect 4219 34790 4265 34842
rect 4265 34790 4275 34842
rect 4299 34790 4329 34842
rect 4329 34790 4341 34842
rect 4341 34790 4355 34842
rect 4379 34790 4393 34842
rect 4393 34790 4405 34842
rect 4405 34790 4435 34842
rect 4459 34790 4469 34842
rect 4469 34790 4515 34842
rect 4219 34788 4275 34790
rect 4299 34788 4355 34790
rect 4379 34788 4435 34790
rect 4459 34788 4515 34790
rect 4219 33754 4275 33756
rect 4299 33754 4355 33756
rect 4379 33754 4435 33756
rect 4459 33754 4515 33756
rect 4219 33702 4265 33754
rect 4265 33702 4275 33754
rect 4299 33702 4329 33754
rect 4329 33702 4341 33754
rect 4341 33702 4355 33754
rect 4379 33702 4393 33754
rect 4393 33702 4405 33754
rect 4405 33702 4435 33754
rect 4459 33702 4469 33754
rect 4469 33702 4515 33754
rect 4219 33700 4275 33702
rect 4299 33700 4355 33702
rect 4379 33700 4435 33702
rect 4459 33700 4515 33702
rect 4219 32666 4275 32668
rect 4299 32666 4355 32668
rect 4379 32666 4435 32668
rect 4459 32666 4515 32668
rect 4219 32614 4265 32666
rect 4265 32614 4275 32666
rect 4299 32614 4329 32666
rect 4329 32614 4341 32666
rect 4341 32614 4355 32666
rect 4379 32614 4393 32666
rect 4393 32614 4405 32666
rect 4405 32614 4435 32666
rect 4459 32614 4469 32666
rect 4469 32614 4515 32666
rect 4219 32612 4275 32614
rect 4299 32612 4355 32614
rect 4379 32612 4435 32614
rect 4459 32612 4515 32614
rect 4219 31578 4275 31580
rect 4299 31578 4355 31580
rect 4379 31578 4435 31580
rect 4459 31578 4515 31580
rect 4219 31526 4265 31578
rect 4265 31526 4275 31578
rect 4299 31526 4329 31578
rect 4329 31526 4341 31578
rect 4341 31526 4355 31578
rect 4379 31526 4393 31578
rect 4393 31526 4405 31578
rect 4405 31526 4435 31578
rect 4459 31526 4469 31578
rect 4469 31526 4515 31578
rect 4219 31524 4275 31526
rect 4299 31524 4355 31526
rect 4379 31524 4435 31526
rect 4459 31524 4515 31526
rect 4219 30490 4275 30492
rect 4299 30490 4355 30492
rect 4379 30490 4435 30492
rect 4459 30490 4515 30492
rect 4219 30438 4265 30490
rect 4265 30438 4275 30490
rect 4299 30438 4329 30490
rect 4329 30438 4341 30490
rect 4341 30438 4355 30490
rect 4379 30438 4393 30490
rect 4393 30438 4405 30490
rect 4405 30438 4435 30490
rect 4459 30438 4469 30490
rect 4469 30438 4515 30490
rect 4219 30436 4275 30438
rect 4299 30436 4355 30438
rect 4379 30436 4435 30438
rect 4459 30436 4515 30438
rect 4219 29402 4275 29404
rect 4299 29402 4355 29404
rect 4379 29402 4435 29404
rect 4459 29402 4515 29404
rect 4219 29350 4265 29402
rect 4265 29350 4275 29402
rect 4299 29350 4329 29402
rect 4329 29350 4341 29402
rect 4341 29350 4355 29402
rect 4379 29350 4393 29402
rect 4393 29350 4405 29402
rect 4405 29350 4435 29402
rect 4459 29350 4469 29402
rect 4469 29350 4515 29402
rect 4219 29348 4275 29350
rect 4299 29348 4355 29350
rect 4379 29348 4435 29350
rect 4459 29348 4515 29350
rect 4219 28314 4275 28316
rect 4299 28314 4355 28316
rect 4379 28314 4435 28316
rect 4459 28314 4515 28316
rect 4219 28262 4265 28314
rect 4265 28262 4275 28314
rect 4299 28262 4329 28314
rect 4329 28262 4341 28314
rect 4341 28262 4355 28314
rect 4379 28262 4393 28314
rect 4393 28262 4405 28314
rect 4405 28262 4435 28314
rect 4459 28262 4469 28314
rect 4469 28262 4515 28314
rect 4219 28260 4275 28262
rect 4299 28260 4355 28262
rect 4379 28260 4435 28262
rect 4459 28260 4515 28262
rect 4219 27226 4275 27228
rect 4299 27226 4355 27228
rect 4379 27226 4435 27228
rect 4459 27226 4515 27228
rect 4219 27174 4265 27226
rect 4265 27174 4275 27226
rect 4299 27174 4329 27226
rect 4329 27174 4341 27226
rect 4341 27174 4355 27226
rect 4379 27174 4393 27226
rect 4393 27174 4405 27226
rect 4405 27174 4435 27226
rect 4459 27174 4469 27226
rect 4469 27174 4515 27226
rect 4219 27172 4275 27174
rect 4299 27172 4355 27174
rect 4379 27172 4435 27174
rect 4459 27172 4515 27174
rect 2588 22330 2644 22332
rect 2668 22330 2724 22332
rect 2748 22330 2804 22332
rect 2828 22330 2884 22332
rect 2588 22278 2634 22330
rect 2634 22278 2644 22330
rect 2668 22278 2698 22330
rect 2698 22278 2710 22330
rect 2710 22278 2724 22330
rect 2748 22278 2762 22330
rect 2762 22278 2774 22330
rect 2774 22278 2804 22330
rect 2828 22278 2838 22330
rect 2838 22278 2884 22330
rect 2588 22276 2644 22278
rect 2668 22276 2724 22278
rect 2748 22276 2804 22278
rect 2828 22276 2884 22278
rect 2042 21664 2098 21720
rect 1582 20712 1638 20768
rect 1490 19488 1546 19544
rect 1398 18944 1454 19000
rect 1398 17312 1454 17368
rect 1674 19896 1730 19952
rect 2870 21392 2926 21448
rect 2588 21242 2644 21244
rect 2668 21242 2724 21244
rect 2748 21242 2804 21244
rect 2828 21242 2884 21244
rect 2588 21190 2634 21242
rect 2634 21190 2644 21242
rect 2668 21190 2698 21242
rect 2698 21190 2710 21242
rect 2710 21190 2724 21242
rect 2748 21190 2762 21242
rect 2762 21190 2774 21242
rect 2774 21190 2804 21242
rect 2828 21190 2838 21242
rect 2838 21190 2884 21242
rect 2588 21188 2644 21190
rect 2668 21188 2724 21190
rect 2748 21188 2804 21190
rect 2828 21188 2884 21190
rect 2588 20154 2644 20156
rect 2668 20154 2724 20156
rect 2748 20154 2804 20156
rect 2828 20154 2884 20156
rect 2588 20102 2634 20154
rect 2634 20102 2644 20154
rect 2668 20102 2698 20154
rect 2698 20102 2710 20154
rect 2710 20102 2724 20154
rect 2748 20102 2762 20154
rect 2762 20102 2774 20154
rect 2774 20102 2804 20154
rect 2828 20102 2838 20154
rect 2838 20102 2884 20154
rect 2588 20100 2644 20102
rect 2668 20100 2724 20102
rect 2748 20100 2804 20102
rect 2828 20100 2884 20102
rect 2588 19066 2644 19068
rect 2668 19066 2724 19068
rect 2748 19066 2804 19068
rect 2828 19066 2884 19068
rect 2588 19014 2634 19066
rect 2634 19014 2644 19066
rect 2668 19014 2698 19066
rect 2698 19014 2710 19066
rect 2710 19014 2724 19066
rect 2748 19014 2762 19066
rect 2762 19014 2774 19066
rect 2774 19014 2804 19066
rect 2828 19014 2838 19066
rect 2838 19014 2884 19066
rect 2588 19012 2644 19014
rect 2668 19012 2724 19014
rect 2748 19012 2804 19014
rect 2828 19012 2884 19014
rect 2588 17978 2644 17980
rect 2668 17978 2724 17980
rect 2748 17978 2804 17980
rect 2828 17978 2884 17980
rect 2588 17926 2634 17978
rect 2634 17926 2644 17978
rect 2668 17926 2698 17978
rect 2698 17926 2710 17978
rect 2710 17926 2724 17978
rect 2748 17926 2762 17978
rect 2762 17926 2774 17978
rect 2774 17926 2804 17978
rect 2828 17926 2838 17978
rect 2838 17926 2884 17978
rect 2588 17924 2644 17926
rect 2668 17924 2724 17926
rect 2748 17924 2804 17926
rect 2828 17924 2884 17926
rect 2870 17620 2872 17640
rect 2872 17620 2924 17640
rect 2924 17620 2926 17640
rect 2870 17584 2926 17620
rect 1398 16224 1454 16280
rect 1490 15000 1546 15056
rect 1398 14456 1454 14512
rect 2588 16890 2644 16892
rect 2668 16890 2724 16892
rect 2748 16890 2804 16892
rect 2828 16890 2884 16892
rect 2588 16838 2634 16890
rect 2634 16838 2644 16890
rect 2668 16838 2698 16890
rect 2698 16838 2710 16890
rect 2710 16838 2724 16890
rect 2748 16838 2762 16890
rect 2762 16838 2774 16890
rect 2774 16838 2804 16890
rect 2828 16838 2838 16890
rect 2838 16838 2884 16890
rect 2588 16836 2644 16838
rect 2668 16836 2724 16838
rect 2748 16836 2804 16838
rect 2828 16836 2884 16838
rect 2226 15816 2282 15872
rect 2588 15802 2644 15804
rect 2668 15802 2724 15804
rect 2748 15802 2804 15804
rect 2828 15802 2884 15804
rect 2588 15750 2634 15802
rect 2634 15750 2644 15802
rect 2668 15750 2698 15802
rect 2698 15750 2710 15802
rect 2710 15750 2724 15802
rect 2748 15750 2762 15802
rect 2762 15750 2774 15802
rect 2774 15750 2804 15802
rect 2828 15750 2838 15802
rect 2838 15750 2884 15802
rect 2588 15748 2644 15750
rect 2668 15748 2724 15750
rect 2748 15748 2804 15750
rect 2828 15748 2884 15750
rect 2226 15444 2228 15464
rect 2228 15444 2280 15464
rect 2280 15444 2282 15464
rect 2226 15408 2282 15444
rect 2588 14714 2644 14716
rect 2668 14714 2724 14716
rect 2748 14714 2804 14716
rect 2828 14714 2884 14716
rect 2588 14662 2634 14714
rect 2634 14662 2644 14714
rect 2668 14662 2698 14714
rect 2698 14662 2710 14714
rect 2710 14662 2724 14714
rect 2748 14662 2762 14714
rect 2762 14662 2774 14714
rect 2774 14662 2804 14714
rect 2828 14662 2838 14714
rect 2838 14662 2884 14714
rect 2588 14660 2644 14662
rect 2668 14660 2724 14662
rect 2748 14660 2804 14662
rect 2828 14660 2884 14662
rect 1398 13096 1454 13152
rect 1490 12280 1546 12336
rect 1398 11736 1454 11792
rect 1398 11328 1454 11384
rect 2318 14048 2374 14104
rect 2226 13640 2282 13696
rect 2226 12688 2282 12744
rect 2588 13626 2644 13628
rect 2668 13626 2724 13628
rect 2748 13626 2804 13628
rect 2828 13626 2884 13628
rect 2588 13574 2634 13626
rect 2634 13574 2644 13626
rect 2668 13574 2698 13626
rect 2698 13574 2710 13626
rect 2710 13574 2724 13626
rect 2748 13574 2762 13626
rect 2762 13574 2774 13626
rect 2774 13574 2804 13626
rect 2828 13574 2838 13626
rect 2838 13574 2884 13626
rect 2588 13572 2644 13574
rect 2668 13572 2724 13574
rect 2748 13572 2804 13574
rect 2828 13572 2884 13574
rect 2588 12538 2644 12540
rect 2668 12538 2724 12540
rect 2748 12538 2804 12540
rect 2828 12538 2884 12540
rect 2588 12486 2634 12538
rect 2634 12486 2644 12538
rect 2668 12486 2698 12538
rect 2698 12486 2710 12538
rect 2710 12486 2724 12538
rect 2748 12486 2762 12538
rect 2762 12486 2774 12538
rect 2774 12486 2804 12538
rect 2828 12486 2838 12538
rect 2838 12486 2884 12538
rect 2588 12484 2644 12486
rect 2668 12484 2724 12486
rect 2748 12484 2804 12486
rect 2828 12484 2884 12486
rect 2588 11450 2644 11452
rect 2668 11450 2724 11452
rect 2748 11450 2804 11452
rect 2828 11450 2884 11452
rect 2588 11398 2634 11450
rect 2634 11398 2644 11450
rect 2668 11398 2698 11450
rect 2698 11398 2710 11450
rect 2710 11398 2724 11450
rect 2748 11398 2762 11450
rect 2762 11398 2774 11450
rect 2774 11398 2804 11450
rect 2828 11398 2838 11450
rect 2838 11398 2884 11450
rect 2588 11396 2644 11398
rect 2668 11396 2724 11398
rect 2748 11396 2804 11398
rect 2828 11396 2884 11398
rect 2588 10362 2644 10364
rect 2668 10362 2724 10364
rect 2748 10362 2804 10364
rect 2828 10362 2884 10364
rect 2588 10310 2634 10362
rect 2634 10310 2644 10362
rect 2668 10310 2698 10362
rect 2698 10310 2710 10362
rect 2710 10310 2724 10362
rect 2748 10310 2762 10362
rect 2762 10310 2774 10362
rect 2774 10310 2804 10362
rect 2828 10310 2838 10362
rect 2838 10310 2884 10362
rect 2588 10308 2644 10310
rect 2668 10308 2724 10310
rect 2748 10308 2804 10310
rect 2828 10308 2884 10310
rect 2588 9274 2644 9276
rect 2668 9274 2724 9276
rect 2748 9274 2804 9276
rect 2828 9274 2884 9276
rect 2588 9222 2634 9274
rect 2634 9222 2644 9274
rect 2668 9222 2698 9274
rect 2698 9222 2710 9274
rect 2710 9222 2724 9274
rect 2748 9222 2762 9274
rect 2762 9222 2774 9274
rect 2774 9222 2804 9274
rect 2828 9222 2838 9274
rect 2838 9222 2884 9274
rect 2588 9220 2644 9222
rect 2668 9220 2724 9222
rect 2748 9220 2804 9222
rect 2828 9220 2884 9222
rect 2588 8186 2644 8188
rect 2668 8186 2724 8188
rect 2748 8186 2804 8188
rect 2828 8186 2884 8188
rect 2588 8134 2634 8186
rect 2634 8134 2644 8186
rect 2668 8134 2698 8186
rect 2698 8134 2710 8186
rect 2710 8134 2724 8186
rect 2748 8134 2762 8186
rect 2762 8134 2774 8186
rect 2774 8134 2804 8186
rect 2828 8134 2838 8186
rect 2838 8134 2884 8186
rect 2588 8132 2644 8134
rect 2668 8132 2724 8134
rect 2748 8132 2804 8134
rect 2828 8132 2884 8134
rect 2588 7098 2644 7100
rect 2668 7098 2724 7100
rect 2748 7098 2804 7100
rect 2828 7098 2884 7100
rect 2588 7046 2634 7098
rect 2634 7046 2644 7098
rect 2668 7046 2698 7098
rect 2698 7046 2710 7098
rect 2710 7046 2724 7098
rect 2748 7046 2762 7098
rect 2762 7046 2774 7098
rect 2774 7046 2804 7098
rect 2828 7046 2838 7098
rect 2838 7046 2884 7098
rect 2588 7044 2644 7046
rect 2668 7044 2724 7046
rect 2748 7044 2804 7046
rect 2828 7044 2884 7046
rect 3330 22072 3386 22128
rect 3790 22616 3846 22672
rect 3514 20304 3570 20360
rect 4219 26138 4275 26140
rect 4299 26138 4355 26140
rect 4379 26138 4435 26140
rect 4459 26138 4515 26140
rect 4219 26086 4265 26138
rect 4265 26086 4275 26138
rect 4299 26086 4329 26138
rect 4329 26086 4341 26138
rect 4341 26086 4355 26138
rect 4379 26086 4393 26138
rect 4393 26086 4405 26138
rect 4405 26086 4435 26138
rect 4459 26086 4469 26138
rect 4469 26086 4515 26138
rect 4219 26084 4275 26086
rect 4299 26084 4355 26086
rect 4379 26084 4435 26086
rect 4459 26084 4515 26086
rect 4219 25050 4275 25052
rect 4299 25050 4355 25052
rect 4379 25050 4435 25052
rect 4459 25050 4515 25052
rect 4219 24998 4265 25050
rect 4265 24998 4275 25050
rect 4299 24998 4329 25050
rect 4329 24998 4341 25050
rect 4341 24998 4355 25050
rect 4379 24998 4393 25050
rect 4393 24998 4405 25050
rect 4405 24998 4435 25050
rect 4459 24998 4469 25050
rect 4469 24998 4515 25050
rect 4219 24996 4275 24998
rect 4299 24996 4355 24998
rect 4379 24996 4435 24998
rect 4459 24996 4515 24998
rect 4802 51584 4858 51640
rect 4986 51176 5042 51232
rect 4894 50904 4950 50960
rect 5851 74554 5907 74556
rect 5931 74554 5987 74556
rect 6011 74554 6067 74556
rect 6091 74554 6147 74556
rect 5851 74502 5897 74554
rect 5897 74502 5907 74554
rect 5931 74502 5961 74554
rect 5961 74502 5973 74554
rect 5973 74502 5987 74554
rect 6011 74502 6025 74554
rect 6025 74502 6037 74554
rect 6037 74502 6067 74554
rect 6091 74502 6101 74554
rect 6101 74502 6147 74554
rect 5851 74500 5907 74502
rect 5931 74500 5987 74502
rect 6011 74500 6067 74502
rect 6091 74500 6147 74502
rect 9115 74554 9171 74556
rect 9195 74554 9251 74556
rect 9275 74554 9331 74556
rect 9355 74554 9411 74556
rect 9115 74502 9161 74554
rect 9161 74502 9171 74554
rect 9195 74502 9225 74554
rect 9225 74502 9237 74554
rect 9237 74502 9251 74554
rect 9275 74502 9289 74554
rect 9289 74502 9301 74554
rect 9301 74502 9331 74554
rect 9355 74502 9365 74554
rect 9365 74502 9411 74554
rect 9115 74500 9171 74502
rect 9195 74500 9251 74502
rect 9275 74500 9331 74502
rect 9355 74500 9411 74502
rect 7483 74010 7539 74012
rect 7563 74010 7619 74012
rect 7643 74010 7699 74012
rect 7723 74010 7779 74012
rect 7483 73958 7529 74010
rect 7529 73958 7539 74010
rect 7563 73958 7593 74010
rect 7593 73958 7605 74010
rect 7605 73958 7619 74010
rect 7643 73958 7657 74010
rect 7657 73958 7669 74010
rect 7669 73958 7699 74010
rect 7723 73958 7733 74010
rect 7733 73958 7779 74010
rect 7483 73956 7539 73958
rect 7563 73956 7619 73958
rect 7643 73956 7699 73958
rect 7723 73956 7779 73958
rect 5851 73466 5907 73468
rect 5931 73466 5987 73468
rect 6011 73466 6067 73468
rect 6091 73466 6147 73468
rect 5851 73414 5897 73466
rect 5897 73414 5907 73466
rect 5931 73414 5961 73466
rect 5961 73414 5973 73466
rect 5973 73414 5987 73466
rect 6011 73414 6025 73466
rect 6025 73414 6037 73466
rect 6037 73414 6067 73466
rect 6091 73414 6101 73466
rect 6101 73414 6147 73466
rect 5851 73412 5907 73414
rect 5931 73412 5987 73414
rect 6011 73412 6067 73414
rect 6091 73412 6147 73414
rect 5446 53624 5502 53680
rect 5354 53080 5410 53136
rect 5354 51312 5410 51368
rect 7483 72922 7539 72924
rect 7563 72922 7619 72924
rect 7643 72922 7699 72924
rect 7723 72922 7779 72924
rect 7483 72870 7529 72922
rect 7529 72870 7539 72922
rect 7563 72870 7593 72922
rect 7593 72870 7605 72922
rect 7605 72870 7619 72922
rect 7643 72870 7657 72922
rect 7657 72870 7669 72922
rect 7669 72870 7699 72922
rect 7723 72870 7733 72922
rect 7733 72870 7779 72922
rect 7483 72868 7539 72870
rect 7563 72868 7619 72870
rect 7643 72868 7699 72870
rect 7723 72868 7779 72870
rect 5851 72378 5907 72380
rect 5931 72378 5987 72380
rect 6011 72378 6067 72380
rect 6091 72378 6147 72380
rect 5851 72326 5897 72378
rect 5897 72326 5907 72378
rect 5931 72326 5961 72378
rect 5961 72326 5973 72378
rect 5973 72326 5987 72378
rect 6011 72326 6025 72378
rect 6025 72326 6037 72378
rect 6037 72326 6067 72378
rect 6091 72326 6101 72378
rect 6101 72326 6147 72378
rect 5851 72324 5907 72326
rect 5931 72324 5987 72326
rect 6011 72324 6067 72326
rect 6091 72324 6147 72326
rect 7483 71834 7539 71836
rect 7563 71834 7619 71836
rect 7643 71834 7699 71836
rect 7723 71834 7779 71836
rect 7483 71782 7529 71834
rect 7529 71782 7539 71834
rect 7563 71782 7593 71834
rect 7593 71782 7605 71834
rect 7605 71782 7619 71834
rect 7643 71782 7657 71834
rect 7657 71782 7669 71834
rect 7669 71782 7699 71834
rect 7723 71782 7733 71834
rect 7733 71782 7779 71834
rect 7483 71780 7539 71782
rect 7563 71780 7619 71782
rect 7643 71780 7699 71782
rect 7723 71780 7779 71782
rect 5851 71290 5907 71292
rect 5931 71290 5987 71292
rect 6011 71290 6067 71292
rect 6091 71290 6147 71292
rect 5851 71238 5897 71290
rect 5897 71238 5907 71290
rect 5931 71238 5961 71290
rect 5961 71238 5973 71290
rect 5973 71238 5987 71290
rect 6011 71238 6025 71290
rect 6025 71238 6037 71290
rect 6037 71238 6067 71290
rect 6091 71238 6101 71290
rect 6101 71238 6147 71290
rect 5851 71236 5907 71238
rect 5931 71236 5987 71238
rect 6011 71236 6067 71238
rect 6091 71236 6147 71238
rect 7483 70746 7539 70748
rect 7563 70746 7619 70748
rect 7643 70746 7699 70748
rect 7723 70746 7779 70748
rect 7483 70694 7529 70746
rect 7529 70694 7539 70746
rect 7563 70694 7593 70746
rect 7593 70694 7605 70746
rect 7605 70694 7619 70746
rect 7643 70694 7657 70746
rect 7657 70694 7669 70746
rect 7669 70694 7699 70746
rect 7723 70694 7733 70746
rect 7733 70694 7779 70746
rect 7483 70692 7539 70694
rect 7563 70692 7619 70694
rect 7643 70692 7699 70694
rect 7723 70692 7779 70694
rect 5851 70202 5907 70204
rect 5931 70202 5987 70204
rect 6011 70202 6067 70204
rect 6091 70202 6147 70204
rect 5851 70150 5897 70202
rect 5897 70150 5907 70202
rect 5931 70150 5961 70202
rect 5961 70150 5973 70202
rect 5973 70150 5987 70202
rect 6011 70150 6025 70202
rect 6025 70150 6037 70202
rect 6037 70150 6067 70202
rect 6091 70150 6101 70202
rect 6101 70150 6147 70202
rect 5851 70148 5907 70150
rect 5931 70148 5987 70150
rect 6011 70148 6067 70150
rect 6091 70148 6147 70150
rect 7483 69658 7539 69660
rect 7563 69658 7619 69660
rect 7643 69658 7699 69660
rect 7723 69658 7779 69660
rect 7483 69606 7529 69658
rect 7529 69606 7539 69658
rect 7563 69606 7593 69658
rect 7593 69606 7605 69658
rect 7605 69606 7619 69658
rect 7643 69606 7657 69658
rect 7657 69606 7669 69658
rect 7669 69606 7699 69658
rect 7723 69606 7733 69658
rect 7733 69606 7779 69658
rect 7483 69604 7539 69606
rect 7563 69604 7619 69606
rect 7643 69604 7699 69606
rect 7723 69604 7779 69606
rect 5851 69114 5907 69116
rect 5931 69114 5987 69116
rect 6011 69114 6067 69116
rect 6091 69114 6147 69116
rect 5851 69062 5897 69114
rect 5897 69062 5907 69114
rect 5931 69062 5961 69114
rect 5961 69062 5973 69114
rect 5973 69062 5987 69114
rect 6011 69062 6025 69114
rect 6025 69062 6037 69114
rect 6037 69062 6067 69114
rect 6091 69062 6101 69114
rect 6101 69062 6147 69114
rect 5851 69060 5907 69062
rect 5931 69060 5987 69062
rect 6011 69060 6067 69062
rect 6091 69060 6147 69062
rect 7483 68570 7539 68572
rect 7563 68570 7619 68572
rect 7643 68570 7699 68572
rect 7723 68570 7779 68572
rect 7483 68518 7529 68570
rect 7529 68518 7539 68570
rect 7563 68518 7593 68570
rect 7593 68518 7605 68570
rect 7605 68518 7619 68570
rect 7643 68518 7657 68570
rect 7657 68518 7669 68570
rect 7669 68518 7699 68570
rect 7723 68518 7733 68570
rect 7733 68518 7779 68570
rect 7483 68516 7539 68518
rect 7563 68516 7619 68518
rect 7643 68516 7699 68518
rect 7723 68516 7779 68518
rect 5851 68026 5907 68028
rect 5931 68026 5987 68028
rect 6011 68026 6067 68028
rect 6091 68026 6147 68028
rect 5851 67974 5897 68026
rect 5897 67974 5907 68026
rect 5931 67974 5961 68026
rect 5961 67974 5973 68026
rect 5973 67974 5987 68026
rect 6011 67974 6025 68026
rect 6025 67974 6037 68026
rect 6037 67974 6067 68026
rect 6091 67974 6101 68026
rect 6101 67974 6147 68026
rect 5851 67972 5907 67974
rect 5931 67972 5987 67974
rect 6011 67972 6067 67974
rect 6091 67972 6147 67974
rect 5851 66938 5907 66940
rect 5931 66938 5987 66940
rect 6011 66938 6067 66940
rect 6091 66938 6147 66940
rect 5851 66886 5897 66938
rect 5897 66886 5907 66938
rect 5931 66886 5961 66938
rect 5961 66886 5973 66938
rect 5973 66886 5987 66938
rect 6011 66886 6025 66938
rect 6025 66886 6037 66938
rect 6037 66886 6067 66938
rect 6091 66886 6101 66938
rect 6101 66886 6147 66938
rect 5851 66884 5907 66886
rect 5931 66884 5987 66886
rect 6011 66884 6067 66886
rect 6091 66884 6147 66886
rect 5851 65850 5907 65852
rect 5931 65850 5987 65852
rect 6011 65850 6067 65852
rect 6091 65850 6147 65852
rect 5851 65798 5897 65850
rect 5897 65798 5907 65850
rect 5931 65798 5961 65850
rect 5961 65798 5973 65850
rect 5973 65798 5987 65850
rect 6011 65798 6025 65850
rect 6025 65798 6037 65850
rect 6037 65798 6067 65850
rect 6091 65798 6101 65850
rect 6101 65798 6147 65850
rect 5851 65796 5907 65798
rect 5931 65796 5987 65798
rect 6011 65796 6067 65798
rect 6091 65796 6147 65798
rect 5851 64762 5907 64764
rect 5931 64762 5987 64764
rect 6011 64762 6067 64764
rect 6091 64762 6147 64764
rect 5851 64710 5897 64762
rect 5897 64710 5907 64762
rect 5931 64710 5961 64762
rect 5961 64710 5973 64762
rect 5973 64710 5987 64762
rect 6011 64710 6025 64762
rect 6025 64710 6037 64762
rect 6037 64710 6067 64762
rect 6091 64710 6101 64762
rect 6101 64710 6147 64762
rect 5851 64708 5907 64710
rect 5931 64708 5987 64710
rect 6011 64708 6067 64710
rect 6091 64708 6147 64710
rect 5851 63674 5907 63676
rect 5931 63674 5987 63676
rect 6011 63674 6067 63676
rect 6091 63674 6147 63676
rect 5851 63622 5897 63674
rect 5897 63622 5907 63674
rect 5931 63622 5961 63674
rect 5961 63622 5973 63674
rect 5973 63622 5987 63674
rect 6011 63622 6025 63674
rect 6025 63622 6037 63674
rect 6037 63622 6067 63674
rect 6091 63622 6101 63674
rect 6101 63622 6147 63674
rect 5851 63620 5907 63622
rect 5931 63620 5987 63622
rect 6011 63620 6067 63622
rect 6091 63620 6147 63622
rect 4219 23962 4275 23964
rect 4299 23962 4355 23964
rect 4379 23962 4435 23964
rect 4459 23962 4515 23964
rect 4219 23910 4265 23962
rect 4265 23910 4275 23962
rect 4299 23910 4329 23962
rect 4329 23910 4341 23962
rect 4341 23910 4355 23962
rect 4379 23910 4393 23962
rect 4393 23910 4405 23962
rect 4405 23910 4435 23962
rect 4459 23910 4469 23962
rect 4469 23910 4515 23962
rect 4219 23908 4275 23910
rect 4299 23908 4355 23910
rect 4379 23908 4435 23910
rect 4459 23908 4515 23910
rect 4219 22874 4275 22876
rect 4299 22874 4355 22876
rect 4379 22874 4435 22876
rect 4459 22874 4515 22876
rect 4219 22822 4265 22874
rect 4265 22822 4275 22874
rect 4299 22822 4329 22874
rect 4329 22822 4341 22874
rect 4341 22822 4355 22874
rect 4379 22822 4393 22874
rect 4393 22822 4405 22874
rect 4405 22822 4435 22874
rect 4459 22822 4469 22874
rect 4469 22822 4515 22874
rect 4219 22820 4275 22822
rect 4299 22820 4355 22822
rect 4379 22820 4435 22822
rect 4459 22820 4515 22822
rect 4219 21786 4275 21788
rect 4299 21786 4355 21788
rect 4379 21786 4435 21788
rect 4459 21786 4515 21788
rect 4219 21734 4265 21786
rect 4265 21734 4275 21786
rect 4299 21734 4329 21786
rect 4329 21734 4341 21786
rect 4341 21734 4355 21786
rect 4379 21734 4393 21786
rect 4393 21734 4405 21786
rect 4405 21734 4435 21786
rect 4459 21734 4469 21786
rect 4469 21734 4515 21786
rect 4219 21732 4275 21734
rect 4299 21732 4355 21734
rect 4379 21732 4435 21734
rect 4459 21732 4515 21734
rect 4219 20698 4275 20700
rect 4299 20698 4355 20700
rect 4379 20698 4435 20700
rect 4459 20698 4515 20700
rect 4219 20646 4265 20698
rect 4265 20646 4275 20698
rect 4299 20646 4329 20698
rect 4329 20646 4341 20698
rect 4341 20646 4355 20698
rect 4379 20646 4393 20698
rect 4393 20646 4405 20698
rect 4405 20646 4435 20698
rect 4459 20646 4469 20698
rect 4469 20646 4515 20698
rect 4219 20644 4275 20646
rect 4299 20644 4355 20646
rect 4379 20644 4435 20646
rect 4459 20644 4515 20646
rect 4219 19610 4275 19612
rect 4299 19610 4355 19612
rect 4379 19610 4435 19612
rect 4459 19610 4515 19612
rect 4219 19558 4265 19610
rect 4265 19558 4275 19610
rect 4299 19558 4329 19610
rect 4329 19558 4341 19610
rect 4341 19558 4355 19610
rect 4379 19558 4393 19610
rect 4393 19558 4405 19610
rect 4405 19558 4435 19610
rect 4459 19558 4469 19610
rect 4469 19558 4515 19610
rect 4219 19556 4275 19558
rect 4299 19556 4355 19558
rect 4379 19556 4435 19558
rect 4459 19556 4515 19558
rect 3514 18128 3570 18184
rect 3974 18536 4030 18592
rect 4219 18522 4275 18524
rect 4299 18522 4355 18524
rect 4379 18522 4435 18524
rect 4459 18522 4515 18524
rect 4219 18470 4265 18522
rect 4265 18470 4275 18522
rect 4299 18470 4329 18522
rect 4329 18470 4341 18522
rect 4341 18470 4355 18522
rect 4379 18470 4393 18522
rect 4393 18470 4405 18522
rect 4405 18470 4435 18522
rect 4459 18470 4469 18522
rect 4469 18470 4515 18522
rect 4219 18468 4275 18470
rect 4299 18468 4355 18470
rect 4379 18468 4435 18470
rect 4459 18468 4515 18470
rect 4219 17434 4275 17436
rect 4299 17434 4355 17436
rect 4379 17434 4435 17436
rect 4459 17434 4515 17436
rect 4219 17382 4265 17434
rect 4265 17382 4275 17434
rect 4299 17382 4329 17434
rect 4329 17382 4341 17434
rect 4341 17382 4355 17434
rect 4379 17382 4393 17434
rect 4393 17382 4405 17434
rect 4405 17382 4435 17434
rect 4459 17382 4469 17434
rect 4469 17382 4515 17434
rect 4219 17380 4275 17382
rect 4299 17380 4355 17382
rect 4379 17380 4435 17382
rect 4459 17380 4515 17382
rect 4219 16346 4275 16348
rect 4299 16346 4355 16348
rect 4379 16346 4435 16348
rect 4459 16346 4515 16348
rect 4219 16294 4265 16346
rect 4265 16294 4275 16346
rect 4299 16294 4329 16346
rect 4329 16294 4341 16346
rect 4341 16294 4355 16346
rect 4379 16294 4393 16346
rect 4393 16294 4405 16346
rect 4405 16294 4435 16346
rect 4459 16294 4469 16346
rect 4469 16294 4515 16346
rect 4219 16292 4275 16294
rect 4299 16292 4355 16294
rect 4379 16292 4435 16294
rect 4459 16292 4515 16294
rect 4219 15258 4275 15260
rect 4299 15258 4355 15260
rect 4379 15258 4435 15260
rect 4459 15258 4515 15260
rect 4219 15206 4265 15258
rect 4265 15206 4275 15258
rect 4299 15206 4329 15258
rect 4329 15206 4341 15258
rect 4341 15206 4355 15258
rect 4379 15206 4393 15258
rect 4393 15206 4405 15258
rect 4405 15206 4435 15258
rect 4459 15206 4469 15258
rect 4469 15206 4515 15258
rect 4219 15204 4275 15206
rect 4299 15204 4355 15206
rect 4379 15204 4435 15206
rect 4459 15204 4515 15206
rect 4219 14170 4275 14172
rect 4299 14170 4355 14172
rect 4379 14170 4435 14172
rect 4459 14170 4515 14172
rect 4219 14118 4265 14170
rect 4265 14118 4275 14170
rect 4299 14118 4329 14170
rect 4329 14118 4341 14170
rect 4341 14118 4355 14170
rect 4379 14118 4393 14170
rect 4393 14118 4405 14170
rect 4405 14118 4435 14170
rect 4459 14118 4469 14170
rect 4469 14118 4515 14170
rect 4219 14116 4275 14118
rect 4299 14116 4355 14118
rect 4379 14116 4435 14118
rect 4459 14116 4515 14118
rect 4219 13082 4275 13084
rect 4299 13082 4355 13084
rect 4379 13082 4435 13084
rect 4459 13082 4515 13084
rect 4219 13030 4265 13082
rect 4265 13030 4275 13082
rect 4299 13030 4329 13082
rect 4329 13030 4341 13082
rect 4341 13030 4355 13082
rect 4379 13030 4393 13082
rect 4393 13030 4405 13082
rect 4405 13030 4435 13082
rect 4459 13030 4469 13082
rect 4469 13030 4515 13082
rect 4219 13028 4275 13030
rect 4299 13028 4355 13030
rect 4379 13028 4435 13030
rect 4459 13028 4515 13030
rect 4219 11994 4275 11996
rect 4299 11994 4355 11996
rect 4379 11994 4435 11996
rect 4459 11994 4515 11996
rect 4219 11942 4265 11994
rect 4265 11942 4275 11994
rect 4299 11942 4329 11994
rect 4329 11942 4341 11994
rect 4341 11942 4355 11994
rect 4379 11942 4393 11994
rect 4393 11942 4405 11994
rect 4405 11942 4435 11994
rect 4459 11942 4469 11994
rect 4469 11942 4515 11994
rect 4219 11940 4275 11942
rect 4299 11940 4355 11942
rect 4379 11940 4435 11942
rect 4459 11940 4515 11942
rect 4219 10906 4275 10908
rect 4299 10906 4355 10908
rect 4379 10906 4435 10908
rect 4459 10906 4515 10908
rect 4219 10854 4265 10906
rect 4265 10854 4275 10906
rect 4299 10854 4329 10906
rect 4329 10854 4341 10906
rect 4341 10854 4355 10906
rect 4379 10854 4393 10906
rect 4393 10854 4405 10906
rect 4405 10854 4435 10906
rect 4459 10854 4469 10906
rect 4469 10854 4515 10906
rect 4219 10852 4275 10854
rect 4299 10852 4355 10854
rect 4379 10852 4435 10854
rect 4459 10852 4515 10854
rect 5446 51040 5502 51096
rect 5354 50904 5410 50960
rect 5262 41384 5318 41440
rect 5851 62586 5907 62588
rect 5931 62586 5987 62588
rect 6011 62586 6067 62588
rect 6091 62586 6147 62588
rect 5851 62534 5897 62586
rect 5897 62534 5907 62586
rect 5931 62534 5961 62586
rect 5961 62534 5973 62586
rect 5973 62534 5987 62586
rect 6011 62534 6025 62586
rect 6025 62534 6037 62586
rect 6037 62534 6067 62586
rect 6091 62534 6101 62586
rect 6101 62534 6147 62586
rect 5851 62532 5907 62534
rect 5931 62532 5987 62534
rect 6011 62532 6067 62534
rect 6091 62532 6147 62534
rect 5851 61498 5907 61500
rect 5931 61498 5987 61500
rect 6011 61498 6067 61500
rect 6091 61498 6147 61500
rect 5851 61446 5897 61498
rect 5897 61446 5907 61498
rect 5931 61446 5961 61498
rect 5961 61446 5973 61498
rect 5973 61446 5987 61498
rect 6011 61446 6025 61498
rect 6025 61446 6037 61498
rect 6037 61446 6067 61498
rect 6091 61446 6101 61498
rect 6101 61446 6147 61498
rect 5851 61444 5907 61446
rect 5931 61444 5987 61446
rect 6011 61444 6067 61446
rect 6091 61444 6147 61446
rect 5851 60410 5907 60412
rect 5931 60410 5987 60412
rect 6011 60410 6067 60412
rect 6091 60410 6147 60412
rect 5851 60358 5897 60410
rect 5897 60358 5907 60410
rect 5931 60358 5961 60410
rect 5961 60358 5973 60410
rect 5973 60358 5987 60410
rect 6011 60358 6025 60410
rect 6025 60358 6037 60410
rect 6037 60358 6067 60410
rect 6091 60358 6101 60410
rect 6101 60358 6147 60410
rect 5851 60356 5907 60358
rect 5931 60356 5987 60358
rect 6011 60356 6067 60358
rect 6091 60356 6147 60358
rect 5851 59322 5907 59324
rect 5931 59322 5987 59324
rect 6011 59322 6067 59324
rect 6091 59322 6147 59324
rect 5851 59270 5897 59322
rect 5897 59270 5907 59322
rect 5931 59270 5961 59322
rect 5961 59270 5973 59322
rect 5973 59270 5987 59322
rect 6011 59270 6025 59322
rect 6025 59270 6037 59322
rect 6037 59270 6067 59322
rect 6091 59270 6101 59322
rect 6101 59270 6147 59322
rect 5851 59268 5907 59270
rect 5931 59268 5987 59270
rect 6011 59268 6067 59270
rect 6091 59268 6147 59270
rect 5851 58234 5907 58236
rect 5931 58234 5987 58236
rect 6011 58234 6067 58236
rect 6091 58234 6147 58236
rect 5851 58182 5897 58234
rect 5897 58182 5907 58234
rect 5931 58182 5961 58234
rect 5961 58182 5973 58234
rect 5973 58182 5987 58234
rect 6011 58182 6025 58234
rect 6025 58182 6037 58234
rect 6037 58182 6067 58234
rect 6091 58182 6101 58234
rect 6101 58182 6147 58234
rect 5851 58180 5907 58182
rect 5931 58180 5987 58182
rect 6011 58180 6067 58182
rect 6091 58180 6147 58182
rect 5851 57146 5907 57148
rect 5931 57146 5987 57148
rect 6011 57146 6067 57148
rect 6091 57146 6147 57148
rect 5851 57094 5897 57146
rect 5897 57094 5907 57146
rect 5931 57094 5961 57146
rect 5961 57094 5973 57146
rect 5973 57094 5987 57146
rect 6011 57094 6025 57146
rect 6025 57094 6037 57146
rect 6037 57094 6067 57146
rect 6091 57094 6101 57146
rect 6101 57094 6147 57146
rect 5851 57092 5907 57094
rect 5931 57092 5987 57094
rect 6011 57092 6067 57094
rect 6091 57092 6147 57094
rect 5851 56058 5907 56060
rect 5931 56058 5987 56060
rect 6011 56058 6067 56060
rect 6091 56058 6147 56060
rect 5851 56006 5897 56058
rect 5897 56006 5907 56058
rect 5931 56006 5961 56058
rect 5961 56006 5973 56058
rect 5973 56006 5987 56058
rect 6011 56006 6025 56058
rect 6025 56006 6037 56058
rect 6037 56006 6067 56058
rect 6091 56006 6101 56058
rect 6101 56006 6147 56058
rect 5851 56004 5907 56006
rect 5931 56004 5987 56006
rect 6011 56004 6067 56006
rect 6091 56004 6147 56006
rect 5851 54970 5907 54972
rect 5931 54970 5987 54972
rect 6011 54970 6067 54972
rect 6091 54970 6147 54972
rect 5851 54918 5897 54970
rect 5897 54918 5907 54970
rect 5931 54918 5961 54970
rect 5961 54918 5973 54970
rect 5973 54918 5987 54970
rect 6011 54918 6025 54970
rect 6025 54918 6037 54970
rect 6037 54918 6067 54970
rect 6091 54918 6101 54970
rect 6101 54918 6147 54970
rect 5851 54916 5907 54918
rect 5931 54916 5987 54918
rect 6011 54916 6067 54918
rect 6091 54916 6147 54918
rect 5851 53882 5907 53884
rect 5931 53882 5987 53884
rect 6011 53882 6067 53884
rect 6091 53882 6147 53884
rect 5851 53830 5897 53882
rect 5897 53830 5907 53882
rect 5931 53830 5961 53882
rect 5961 53830 5973 53882
rect 5973 53830 5987 53882
rect 6011 53830 6025 53882
rect 6025 53830 6037 53882
rect 6037 53830 6067 53882
rect 6091 53830 6101 53882
rect 6101 53830 6147 53882
rect 5851 53828 5907 53830
rect 5931 53828 5987 53830
rect 6011 53828 6067 53830
rect 6091 53828 6147 53830
rect 5851 52794 5907 52796
rect 5931 52794 5987 52796
rect 6011 52794 6067 52796
rect 6091 52794 6147 52796
rect 5851 52742 5897 52794
rect 5897 52742 5907 52794
rect 5931 52742 5961 52794
rect 5961 52742 5973 52794
rect 5973 52742 5987 52794
rect 6011 52742 6025 52794
rect 6025 52742 6037 52794
rect 6037 52742 6067 52794
rect 6091 52742 6101 52794
rect 6101 52742 6147 52794
rect 5851 52740 5907 52742
rect 5931 52740 5987 52742
rect 6011 52740 6067 52742
rect 6091 52740 6147 52742
rect 5851 51706 5907 51708
rect 5931 51706 5987 51708
rect 6011 51706 6067 51708
rect 6091 51706 6147 51708
rect 5851 51654 5897 51706
rect 5897 51654 5907 51706
rect 5931 51654 5961 51706
rect 5961 51654 5973 51706
rect 5973 51654 5987 51706
rect 6011 51654 6025 51706
rect 6025 51654 6037 51706
rect 6037 51654 6067 51706
rect 6091 51654 6101 51706
rect 6101 51654 6147 51706
rect 5851 51652 5907 51654
rect 5931 51652 5987 51654
rect 6011 51652 6067 51654
rect 6091 51652 6147 51654
rect 5851 50618 5907 50620
rect 5931 50618 5987 50620
rect 6011 50618 6067 50620
rect 6091 50618 6147 50620
rect 5851 50566 5897 50618
rect 5897 50566 5907 50618
rect 5931 50566 5961 50618
rect 5961 50566 5973 50618
rect 5973 50566 5987 50618
rect 6011 50566 6025 50618
rect 6025 50566 6037 50618
rect 6037 50566 6067 50618
rect 6091 50566 6101 50618
rect 6101 50566 6147 50618
rect 5851 50564 5907 50566
rect 5931 50564 5987 50566
rect 6011 50564 6067 50566
rect 6091 50564 6147 50566
rect 5851 49530 5907 49532
rect 5931 49530 5987 49532
rect 6011 49530 6067 49532
rect 6091 49530 6147 49532
rect 5851 49478 5897 49530
rect 5897 49478 5907 49530
rect 5931 49478 5961 49530
rect 5961 49478 5973 49530
rect 5973 49478 5987 49530
rect 6011 49478 6025 49530
rect 6025 49478 6037 49530
rect 6037 49478 6067 49530
rect 6091 49478 6101 49530
rect 6101 49478 6147 49530
rect 5851 49476 5907 49478
rect 5931 49476 5987 49478
rect 6011 49476 6067 49478
rect 6091 49476 6147 49478
rect 5851 48442 5907 48444
rect 5931 48442 5987 48444
rect 6011 48442 6067 48444
rect 6091 48442 6147 48444
rect 5851 48390 5897 48442
rect 5897 48390 5907 48442
rect 5931 48390 5961 48442
rect 5961 48390 5973 48442
rect 5973 48390 5987 48442
rect 6011 48390 6025 48442
rect 6025 48390 6037 48442
rect 6037 48390 6067 48442
rect 6091 48390 6101 48442
rect 6101 48390 6147 48442
rect 5851 48388 5907 48390
rect 5931 48388 5987 48390
rect 6011 48388 6067 48390
rect 6091 48388 6147 48390
rect 5851 47354 5907 47356
rect 5931 47354 5987 47356
rect 6011 47354 6067 47356
rect 6091 47354 6147 47356
rect 5851 47302 5897 47354
rect 5897 47302 5907 47354
rect 5931 47302 5961 47354
rect 5961 47302 5973 47354
rect 5973 47302 5987 47354
rect 6011 47302 6025 47354
rect 6025 47302 6037 47354
rect 6037 47302 6067 47354
rect 6091 47302 6101 47354
rect 6101 47302 6147 47354
rect 5851 47300 5907 47302
rect 5931 47300 5987 47302
rect 6011 47300 6067 47302
rect 6091 47300 6147 47302
rect 5851 46266 5907 46268
rect 5931 46266 5987 46268
rect 6011 46266 6067 46268
rect 6091 46266 6147 46268
rect 5851 46214 5897 46266
rect 5897 46214 5907 46266
rect 5931 46214 5961 46266
rect 5961 46214 5973 46266
rect 5973 46214 5987 46266
rect 6011 46214 6025 46266
rect 6025 46214 6037 46266
rect 6037 46214 6067 46266
rect 6091 46214 6101 46266
rect 6101 46214 6147 46266
rect 5851 46212 5907 46214
rect 5931 46212 5987 46214
rect 6011 46212 6067 46214
rect 6091 46212 6147 46214
rect 5851 45178 5907 45180
rect 5931 45178 5987 45180
rect 6011 45178 6067 45180
rect 6091 45178 6147 45180
rect 5851 45126 5897 45178
rect 5897 45126 5907 45178
rect 5931 45126 5961 45178
rect 5961 45126 5973 45178
rect 5973 45126 5987 45178
rect 6011 45126 6025 45178
rect 6025 45126 6037 45178
rect 6037 45126 6067 45178
rect 6091 45126 6101 45178
rect 6101 45126 6147 45178
rect 5851 45124 5907 45126
rect 5931 45124 5987 45126
rect 6011 45124 6067 45126
rect 6091 45124 6147 45126
rect 5851 44090 5907 44092
rect 5931 44090 5987 44092
rect 6011 44090 6067 44092
rect 6091 44090 6147 44092
rect 5851 44038 5897 44090
rect 5897 44038 5907 44090
rect 5931 44038 5961 44090
rect 5961 44038 5973 44090
rect 5973 44038 5987 44090
rect 6011 44038 6025 44090
rect 6025 44038 6037 44090
rect 6037 44038 6067 44090
rect 6091 44038 6101 44090
rect 6101 44038 6147 44090
rect 5851 44036 5907 44038
rect 5931 44036 5987 44038
rect 6011 44036 6067 44038
rect 6091 44036 6147 44038
rect 5851 43002 5907 43004
rect 5931 43002 5987 43004
rect 6011 43002 6067 43004
rect 6091 43002 6147 43004
rect 5851 42950 5897 43002
rect 5897 42950 5907 43002
rect 5931 42950 5961 43002
rect 5961 42950 5973 43002
rect 5973 42950 5987 43002
rect 6011 42950 6025 43002
rect 6025 42950 6037 43002
rect 6037 42950 6067 43002
rect 6091 42950 6101 43002
rect 6101 42950 6147 43002
rect 5851 42948 5907 42950
rect 5931 42948 5987 42950
rect 6011 42948 6067 42950
rect 6091 42948 6147 42950
rect 5851 41914 5907 41916
rect 5931 41914 5987 41916
rect 6011 41914 6067 41916
rect 6091 41914 6147 41916
rect 5851 41862 5897 41914
rect 5897 41862 5907 41914
rect 5931 41862 5961 41914
rect 5961 41862 5973 41914
rect 5973 41862 5987 41914
rect 6011 41862 6025 41914
rect 6025 41862 6037 41914
rect 6037 41862 6067 41914
rect 6091 41862 6101 41914
rect 6101 41862 6147 41914
rect 5851 41860 5907 41862
rect 5931 41860 5987 41862
rect 6011 41860 6067 41862
rect 6091 41860 6147 41862
rect 5851 40826 5907 40828
rect 5931 40826 5987 40828
rect 6011 40826 6067 40828
rect 6091 40826 6147 40828
rect 5851 40774 5897 40826
rect 5897 40774 5907 40826
rect 5931 40774 5961 40826
rect 5961 40774 5973 40826
rect 5973 40774 5987 40826
rect 6011 40774 6025 40826
rect 6025 40774 6037 40826
rect 6037 40774 6067 40826
rect 6091 40774 6101 40826
rect 6101 40774 6147 40826
rect 5851 40772 5907 40774
rect 5931 40772 5987 40774
rect 6011 40772 6067 40774
rect 6091 40772 6147 40774
rect 5851 39738 5907 39740
rect 5931 39738 5987 39740
rect 6011 39738 6067 39740
rect 6091 39738 6147 39740
rect 5851 39686 5897 39738
rect 5897 39686 5907 39738
rect 5931 39686 5961 39738
rect 5961 39686 5973 39738
rect 5973 39686 5987 39738
rect 6011 39686 6025 39738
rect 6025 39686 6037 39738
rect 6037 39686 6067 39738
rect 6091 39686 6101 39738
rect 6101 39686 6147 39738
rect 5851 39684 5907 39686
rect 5931 39684 5987 39686
rect 6011 39684 6067 39686
rect 6091 39684 6147 39686
rect 5851 38650 5907 38652
rect 5931 38650 5987 38652
rect 6011 38650 6067 38652
rect 6091 38650 6147 38652
rect 5851 38598 5897 38650
rect 5897 38598 5907 38650
rect 5931 38598 5961 38650
rect 5961 38598 5973 38650
rect 5973 38598 5987 38650
rect 6011 38598 6025 38650
rect 6025 38598 6037 38650
rect 6037 38598 6067 38650
rect 6091 38598 6101 38650
rect 6101 38598 6147 38650
rect 5851 38596 5907 38598
rect 5931 38596 5987 38598
rect 6011 38596 6067 38598
rect 6091 38596 6147 38598
rect 5851 37562 5907 37564
rect 5931 37562 5987 37564
rect 6011 37562 6067 37564
rect 6091 37562 6147 37564
rect 5851 37510 5897 37562
rect 5897 37510 5907 37562
rect 5931 37510 5961 37562
rect 5961 37510 5973 37562
rect 5973 37510 5987 37562
rect 6011 37510 6025 37562
rect 6025 37510 6037 37562
rect 6037 37510 6067 37562
rect 6091 37510 6101 37562
rect 6101 37510 6147 37562
rect 5851 37508 5907 37510
rect 5931 37508 5987 37510
rect 6011 37508 6067 37510
rect 6091 37508 6147 37510
rect 5851 36474 5907 36476
rect 5931 36474 5987 36476
rect 6011 36474 6067 36476
rect 6091 36474 6147 36476
rect 5851 36422 5897 36474
rect 5897 36422 5907 36474
rect 5931 36422 5961 36474
rect 5961 36422 5973 36474
rect 5973 36422 5987 36474
rect 6011 36422 6025 36474
rect 6025 36422 6037 36474
rect 6037 36422 6067 36474
rect 6091 36422 6101 36474
rect 6101 36422 6147 36474
rect 5851 36420 5907 36422
rect 5931 36420 5987 36422
rect 6011 36420 6067 36422
rect 6091 36420 6147 36422
rect 5851 35386 5907 35388
rect 5931 35386 5987 35388
rect 6011 35386 6067 35388
rect 6091 35386 6147 35388
rect 5851 35334 5897 35386
rect 5897 35334 5907 35386
rect 5931 35334 5961 35386
rect 5961 35334 5973 35386
rect 5973 35334 5987 35386
rect 6011 35334 6025 35386
rect 6025 35334 6037 35386
rect 6037 35334 6067 35386
rect 6091 35334 6101 35386
rect 6101 35334 6147 35386
rect 5851 35332 5907 35334
rect 5931 35332 5987 35334
rect 6011 35332 6067 35334
rect 6091 35332 6147 35334
rect 5851 34298 5907 34300
rect 5931 34298 5987 34300
rect 6011 34298 6067 34300
rect 6091 34298 6147 34300
rect 5851 34246 5897 34298
rect 5897 34246 5907 34298
rect 5931 34246 5961 34298
rect 5961 34246 5973 34298
rect 5973 34246 5987 34298
rect 6011 34246 6025 34298
rect 6025 34246 6037 34298
rect 6037 34246 6067 34298
rect 6091 34246 6101 34298
rect 6101 34246 6147 34298
rect 5851 34244 5907 34246
rect 5931 34244 5987 34246
rect 6011 34244 6067 34246
rect 6091 34244 6147 34246
rect 5851 33210 5907 33212
rect 5931 33210 5987 33212
rect 6011 33210 6067 33212
rect 6091 33210 6147 33212
rect 5851 33158 5897 33210
rect 5897 33158 5907 33210
rect 5931 33158 5961 33210
rect 5961 33158 5973 33210
rect 5973 33158 5987 33210
rect 6011 33158 6025 33210
rect 6025 33158 6037 33210
rect 6037 33158 6067 33210
rect 6091 33158 6101 33210
rect 6101 33158 6147 33210
rect 5851 33156 5907 33158
rect 5931 33156 5987 33158
rect 6011 33156 6067 33158
rect 6091 33156 6147 33158
rect 5851 32122 5907 32124
rect 5931 32122 5987 32124
rect 6011 32122 6067 32124
rect 6091 32122 6147 32124
rect 5851 32070 5897 32122
rect 5897 32070 5907 32122
rect 5931 32070 5961 32122
rect 5961 32070 5973 32122
rect 5973 32070 5987 32122
rect 6011 32070 6025 32122
rect 6025 32070 6037 32122
rect 6037 32070 6067 32122
rect 6091 32070 6101 32122
rect 6101 32070 6147 32122
rect 5851 32068 5907 32070
rect 5931 32068 5987 32070
rect 6011 32068 6067 32070
rect 6091 32068 6147 32070
rect 5851 31034 5907 31036
rect 5931 31034 5987 31036
rect 6011 31034 6067 31036
rect 6091 31034 6147 31036
rect 5851 30982 5897 31034
rect 5897 30982 5907 31034
rect 5931 30982 5961 31034
rect 5961 30982 5973 31034
rect 5973 30982 5987 31034
rect 6011 30982 6025 31034
rect 6025 30982 6037 31034
rect 6037 30982 6067 31034
rect 6091 30982 6101 31034
rect 6101 30982 6147 31034
rect 5851 30980 5907 30982
rect 5931 30980 5987 30982
rect 6011 30980 6067 30982
rect 6091 30980 6147 30982
rect 5851 29946 5907 29948
rect 5931 29946 5987 29948
rect 6011 29946 6067 29948
rect 6091 29946 6147 29948
rect 5851 29894 5897 29946
rect 5897 29894 5907 29946
rect 5931 29894 5961 29946
rect 5961 29894 5973 29946
rect 5973 29894 5987 29946
rect 6011 29894 6025 29946
rect 6025 29894 6037 29946
rect 6037 29894 6067 29946
rect 6091 29894 6101 29946
rect 6101 29894 6147 29946
rect 5851 29892 5907 29894
rect 5931 29892 5987 29894
rect 6011 29892 6067 29894
rect 6091 29892 6147 29894
rect 5851 28858 5907 28860
rect 5931 28858 5987 28860
rect 6011 28858 6067 28860
rect 6091 28858 6147 28860
rect 5851 28806 5897 28858
rect 5897 28806 5907 28858
rect 5931 28806 5961 28858
rect 5961 28806 5973 28858
rect 5973 28806 5987 28858
rect 6011 28806 6025 28858
rect 6025 28806 6037 28858
rect 6037 28806 6067 28858
rect 6091 28806 6101 28858
rect 6101 28806 6147 28858
rect 5851 28804 5907 28806
rect 5931 28804 5987 28806
rect 6011 28804 6067 28806
rect 6091 28804 6147 28806
rect 5851 27770 5907 27772
rect 5931 27770 5987 27772
rect 6011 27770 6067 27772
rect 6091 27770 6147 27772
rect 5851 27718 5897 27770
rect 5897 27718 5907 27770
rect 5931 27718 5961 27770
rect 5961 27718 5973 27770
rect 5973 27718 5987 27770
rect 6011 27718 6025 27770
rect 6025 27718 6037 27770
rect 6037 27718 6067 27770
rect 6091 27718 6101 27770
rect 6101 27718 6147 27770
rect 5851 27716 5907 27718
rect 5931 27716 5987 27718
rect 6011 27716 6067 27718
rect 6091 27716 6147 27718
rect 5851 26682 5907 26684
rect 5931 26682 5987 26684
rect 6011 26682 6067 26684
rect 6091 26682 6147 26684
rect 5851 26630 5897 26682
rect 5897 26630 5907 26682
rect 5931 26630 5961 26682
rect 5961 26630 5973 26682
rect 5973 26630 5987 26682
rect 6011 26630 6025 26682
rect 6025 26630 6037 26682
rect 6037 26630 6067 26682
rect 6091 26630 6101 26682
rect 6101 26630 6147 26682
rect 5851 26628 5907 26630
rect 5931 26628 5987 26630
rect 6011 26628 6067 26630
rect 6091 26628 6147 26630
rect 5851 25594 5907 25596
rect 5931 25594 5987 25596
rect 6011 25594 6067 25596
rect 6091 25594 6147 25596
rect 5851 25542 5897 25594
rect 5897 25542 5907 25594
rect 5931 25542 5961 25594
rect 5961 25542 5973 25594
rect 5973 25542 5987 25594
rect 6011 25542 6025 25594
rect 6025 25542 6037 25594
rect 6037 25542 6067 25594
rect 6091 25542 6101 25594
rect 6101 25542 6147 25594
rect 5851 25540 5907 25542
rect 5931 25540 5987 25542
rect 6011 25540 6067 25542
rect 6091 25540 6147 25542
rect 5851 24506 5907 24508
rect 5931 24506 5987 24508
rect 6011 24506 6067 24508
rect 6091 24506 6147 24508
rect 5851 24454 5897 24506
rect 5897 24454 5907 24506
rect 5931 24454 5961 24506
rect 5961 24454 5973 24506
rect 5973 24454 5987 24506
rect 6011 24454 6025 24506
rect 6025 24454 6037 24506
rect 6037 24454 6067 24506
rect 6091 24454 6101 24506
rect 6101 24454 6147 24506
rect 5851 24452 5907 24454
rect 5931 24452 5987 24454
rect 6011 24452 6067 24454
rect 6091 24452 6147 24454
rect 5851 23418 5907 23420
rect 5931 23418 5987 23420
rect 6011 23418 6067 23420
rect 6091 23418 6147 23420
rect 5851 23366 5897 23418
rect 5897 23366 5907 23418
rect 5931 23366 5961 23418
rect 5961 23366 5973 23418
rect 5973 23366 5987 23418
rect 6011 23366 6025 23418
rect 6025 23366 6037 23418
rect 6037 23366 6067 23418
rect 6091 23366 6101 23418
rect 6101 23366 6147 23418
rect 5851 23364 5907 23366
rect 5931 23364 5987 23366
rect 6011 23364 6067 23366
rect 6091 23364 6147 23366
rect 5851 22330 5907 22332
rect 5931 22330 5987 22332
rect 6011 22330 6067 22332
rect 6091 22330 6147 22332
rect 5851 22278 5897 22330
rect 5897 22278 5907 22330
rect 5931 22278 5961 22330
rect 5961 22278 5973 22330
rect 5973 22278 5987 22330
rect 6011 22278 6025 22330
rect 6025 22278 6037 22330
rect 6037 22278 6067 22330
rect 6091 22278 6101 22330
rect 6101 22278 6147 22330
rect 5851 22276 5907 22278
rect 5931 22276 5987 22278
rect 6011 22276 6067 22278
rect 6091 22276 6147 22278
rect 5851 21242 5907 21244
rect 5931 21242 5987 21244
rect 6011 21242 6067 21244
rect 6091 21242 6147 21244
rect 5851 21190 5897 21242
rect 5897 21190 5907 21242
rect 5931 21190 5961 21242
rect 5961 21190 5973 21242
rect 5973 21190 5987 21242
rect 6011 21190 6025 21242
rect 6025 21190 6037 21242
rect 6037 21190 6067 21242
rect 6091 21190 6101 21242
rect 6101 21190 6147 21242
rect 5851 21188 5907 21190
rect 5931 21188 5987 21190
rect 6011 21188 6067 21190
rect 6091 21188 6147 21190
rect 5851 20154 5907 20156
rect 5931 20154 5987 20156
rect 6011 20154 6067 20156
rect 6091 20154 6147 20156
rect 5851 20102 5897 20154
rect 5897 20102 5907 20154
rect 5931 20102 5961 20154
rect 5961 20102 5973 20154
rect 5973 20102 5987 20154
rect 6011 20102 6025 20154
rect 6025 20102 6037 20154
rect 6037 20102 6067 20154
rect 6091 20102 6101 20154
rect 6101 20102 6147 20154
rect 5851 20100 5907 20102
rect 5931 20100 5987 20102
rect 6011 20100 6067 20102
rect 6091 20100 6147 20102
rect 5851 19066 5907 19068
rect 5931 19066 5987 19068
rect 6011 19066 6067 19068
rect 6091 19066 6147 19068
rect 5851 19014 5897 19066
rect 5897 19014 5907 19066
rect 5931 19014 5961 19066
rect 5961 19014 5973 19066
rect 5973 19014 5987 19066
rect 6011 19014 6025 19066
rect 6025 19014 6037 19066
rect 6037 19014 6067 19066
rect 6091 19014 6101 19066
rect 6101 19014 6147 19066
rect 5851 19012 5907 19014
rect 5931 19012 5987 19014
rect 6011 19012 6067 19014
rect 6091 19012 6147 19014
rect 5851 17978 5907 17980
rect 5931 17978 5987 17980
rect 6011 17978 6067 17980
rect 6091 17978 6147 17980
rect 5851 17926 5897 17978
rect 5897 17926 5907 17978
rect 5931 17926 5961 17978
rect 5961 17926 5973 17978
rect 5973 17926 5987 17978
rect 6011 17926 6025 17978
rect 6025 17926 6037 17978
rect 6037 17926 6067 17978
rect 6091 17926 6101 17978
rect 6101 17926 6147 17978
rect 5851 17924 5907 17926
rect 5931 17924 5987 17926
rect 6011 17924 6067 17926
rect 6091 17924 6147 17926
rect 6826 48728 6882 48784
rect 6734 46280 6790 46336
rect 5851 16890 5907 16892
rect 5931 16890 5987 16892
rect 6011 16890 6067 16892
rect 6091 16890 6147 16892
rect 5851 16838 5897 16890
rect 5897 16838 5907 16890
rect 5931 16838 5961 16890
rect 5961 16838 5973 16890
rect 5973 16838 5987 16890
rect 6011 16838 6025 16890
rect 6025 16838 6037 16890
rect 6037 16838 6067 16890
rect 6091 16838 6101 16890
rect 6101 16838 6147 16890
rect 5851 16836 5907 16838
rect 5931 16836 5987 16838
rect 6011 16836 6067 16838
rect 6091 16836 6147 16838
rect 5851 15802 5907 15804
rect 5931 15802 5987 15804
rect 6011 15802 6067 15804
rect 6091 15802 6147 15804
rect 5851 15750 5897 15802
rect 5897 15750 5907 15802
rect 5931 15750 5961 15802
rect 5961 15750 5973 15802
rect 5973 15750 5987 15802
rect 6011 15750 6025 15802
rect 6025 15750 6037 15802
rect 6037 15750 6067 15802
rect 6091 15750 6101 15802
rect 6101 15750 6147 15802
rect 5851 15748 5907 15750
rect 5931 15748 5987 15750
rect 6011 15748 6067 15750
rect 6091 15748 6147 15750
rect 5851 14714 5907 14716
rect 5931 14714 5987 14716
rect 6011 14714 6067 14716
rect 6091 14714 6147 14716
rect 5851 14662 5897 14714
rect 5897 14662 5907 14714
rect 5931 14662 5961 14714
rect 5961 14662 5973 14714
rect 5973 14662 5987 14714
rect 6011 14662 6025 14714
rect 6025 14662 6037 14714
rect 6037 14662 6067 14714
rect 6091 14662 6101 14714
rect 6101 14662 6147 14714
rect 5851 14660 5907 14662
rect 5931 14660 5987 14662
rect 6011 14660 6067 14662
rect 6091 14660 6147 14662
rect 5851 13626 5907 13628
rect 5931 13626 5987 13628
rect 6011 13626 6067 13628
rect 6091 13626 6147 13628
rect 5851 13574 5897 13626
rect 5897 13574 5907 13626
rect 5931 13574 5961 13626
rect 5961 13574 5973 13626
rect 5973 13574 5987 13626
rect 6011 13574 6025 13626
rect 6025 13574 6037 13626
rect 6037 13574 6067 13626
rect 6091 13574 6101 13626
rect 6101 13574 6147 13626
rect 5851 13572 5907 13574
rect 5931 13572 5987 13574
rect 6011 13572 6067 13574
rect 6091 13572 6147 13574
rect 5851 12538 5907 12540
rect 5931 12538 5987 12540
rect 6011 12538 6067 12540
rect 6091 12538 6147 12540
rect 5851 12486 5897 12538
rect 5897 12486 5907 12538
rect 5931 12486 5961 12538
rect 5961 12486 5973 12538
rect 5973 12486 5987 12538
rect 6011 12486 6025 12538
rect 6025 12486 6037 12538
rect 6037 12486 6067 12538
rect 6091 12486 6101 12538
rect 6101 12486 6147 12538
rect 5851 12484 5907 12486
rect 5931 12484 5987 12486
rect 6011 12484 6067 12486
rect 6091 12484 6147 12486
rect 5851 11450 5907 11452
rect 5931 11450 5987 11452
rect 6011 11450 6067 11452
rect 6091 11450 6147 11452
rect 5851 11398 5897 11450
rect 5897 11398 5907 11450
rect 5931 11398 5961 11450
rect 5961 11398 5973 11450
rect 5973 11398 5987 11450
rect 6011 11398 6025 11450
rect 6025 11398 6037 11450
rect 6037 11398 6067 11450
rect 6091 11398 6101 11450
rect 6101 11398 6147 11450
rect 5851 11396 5907 11398
rect 5931 11396 5987 11398
rect 6011 11396 6067 11398
rect 6091 11396 6147 11398
rect 4219 9818 4275 9820
rect 4299 9818 4355 9820
rect 4379 9818 4435 9820
rect 4459 9818 4515 9820
rect 4219 9766 4265 9818
rect 4265 9766 4275 9818
rect 4299 9766 4329 9818
rect 4329 9766 4341 9818
rect 4341 9766 4355 9818
rect 4379 9766 4393 9818
rect 4393 9766 4405 9818
rect 4405 9766 4435 9818
rect 4459 9766 4469 9818
rect 4469 9766 4515 9818
rect 4219 9764 4275 9766
rect 4299 9764 4355 9766
rect 4379 9764 4435 9766
rect 4459 9764 4515 9766
rect 5851 10362 5907 10364
rect 5931 10362 5987 10364
rect 6011 10362 6067 10364
rect 6091 10362 6147 10364
rect 5851 10310 5897 10362
rect 5897 10310 5907 10362
rect 5931 10310 5961 10362
rect 5961 10310 5973 10362
rect 5973 10310 5987 10362
rect 6011 10310 6025 10362
rect 6025 10310 6037 10362
rect 6037 10310 6067 10362
rect 6091 10310 6101 10362
rect 6101 10310 6147 10362
rect 5851 10308 5907 10310
rect 5931 10308 5987 10310
rect 6011 10308 6067 10310
rect 6091 10308 6147 10310
rect 4219 8730 4275 8732
rect 4299 8730 4355 8732
rect 4379 8730 4435 8732
rect 4459 8730 4515 8732
rect 4219 8678 4265 8730
rect 4265 8678 4275 8730
rect 4299 8678 4329 8730
rect 4329 8678 4341 8730
rect 4341 8678 4355 8730
rect 4379 8678 4393 8730
rect 4393 8678 4405 8730
rect 4405 8678 4435 8730
rect 4459 8678 4469 8730
rect 4469 8678 4515 8730
rect 4219 8676 4275 8678
rect 4299 8676 4355 8678
rect 4379 8676 4435 8678
rect 4459 8676 4515 8678
rect 1398 3712 1454 3768
rect 1214 3304 1270 3360
rect 1306 2760 1362 2816
rect 2588 6010 2644 6012
rect 2668 6010 2724 6012
rect 2748 6010 2804 6012
rect 2828 6010 2884 6012
rect 2588 5958 2634 6010
rect 2634 5958 2644 6010
rect 2668 5958 2698 6010
rect 2698 5958 2710 6010
rect 2710 5958 2724 6010
rect 2748 5958 2762 6010
rect 2762 5958 2774 6010
rect 2774 5958 2804 6010
rect 2828 5958 2838 6010
rect 2838 5958 2884 6010
rect 2588 5956 2644 5958
rect 2668 5956 2724 5958
rect 2748 5956 2804 5958
rect 2828 5956 2884 5958
rect 4219 7642 4275 7644
rect 4299 7642 4355 7644
rect 4379 7642 4435 7644
rect 4459 7642 4515 7644
rect 4219 7590 4265 7642
rect 4265 7590 4275 7642
rect 4299 7590 4329 7642
rect 4329 7590 4341 7642
rect 4341 7590 4355 7642
rect 4379 7590 4393 7642
rect 4393 7590 4405 7642
rect 4405 7590 4435 7642
rect 4459 7590 4469 7642
rect 4469 7590 4515 7642
rect 4219 7588 4275 7590
rect 4299 7588 4355 7590
rect 4379 7588 4435 7590
rect 4459 7588 4515 7590
rect 5851 9274 5907 9276
rect 5931 9274 5987 9276
rect 6011 9274 6067 9276
rect 6091 9274 6147 9276
rect 5851 9222 5897 9274
rect 5897 9222 5907 9274
rect 5931 9222 5961 9274
rect 5961 9222 5973 9274
rect 5973 9222 5987 9274
rect 6011 9222 6025 9274
rect 6025 9222 6037 9274
rect 6037 9222 6067 9274
rect 6091 9222 6101 9274
rect 6101 9222 6147 9274
rect 5851 9220 5907 9222
rect 5931 9220 5987 9222
rect 6011 9220 6067 9222
rect 6091 9220 6147 9222
rect 5851 8186 5907 8188
rect 5931 8186 5987 8188
rect 6011 8186 6067 8188
rect 6091 8186 6147 8188
rect 5851 8134 5897 8186
rect 5897 8134 5907 8186
rect 5931 8134 5961 8186
rect 5961 8134 5973 8186
rect 5973 8134 5987 8186
rect 6011 8134 6025 8186
rect 6025 8134 6037 8186
rect 6037 8134 6067 8186
rect 6091 8134 6101 8186
rect 6101 8134 6147 8186
rect 5851 8132 5907 8134
rect 5931 8132 5987 8134
rect 6011 8132 6067 8134
rect 6091 8132 6147 8134
rect 5851 7098 5907 7100
rect 5931 7098 5987 7100
rect 6011 7098 6067 7100
rect 6091 7098 6147 7100
rect 5851 7046 5897 7098
rect 5897 7046 5907 7098
rect 5931 7046 5961 7098
rect 5961 7046 5973 7098
rect 5973 7046 5987 7098
rect 6011 7046 6025 7098
rect 6025 7046 6037 7098
rect 6037 7046 6067 7098
rect 6091 7046 6101 7098
rect 6101 7046 6147 7098
rect 5851 7044 5907 7046
rect 5931 7044 5987 7046
rect 6011 7044 6067 7046
rect 6091 7044 6147 7046
rect 4219 6554 4275 6556
rect 4299 6554 4355 6556
rect 4379 6554 4435 6556
rect 4459 6554 4515 6556
rect 4219 6502 4265 6554
rect 4265 6502 4275 6554
rect 4299 6502 4329 6554
rect 4329 6502 4341 6554
rect 4341 6502 4355 6554
rect 4379 6502 4393 6554
rect 4393 6502 4405 6554
rect 4405 6502 4435 6554
rect 4459 6502 4469 6554
rect 4469 6502 4515 6554
rect 4219 6500 4275 6502
rect 4299 6500 4355 6502
rect 4379 6500 4435 6502
rect 4459 6500 4515 6502
rect 2588 4922 2644 4924
rect 2668 4922 2724 4924
rect 2748 4922 2804 4924
rect 2828 4922 2884 4924
rect 2588 4870 2634 4922
rect 2634 4870 2644 4922
rect 2668 4870 2698 4922
rect 2698 4870 2710 4922
rect 2710 4870 2724 4922
rect 2748 4870 2762 4922
rect 2762 4870 2774 4922
rect 2774 4870 2804 4922
rect 2828 4870 2838 4922
rect 2838 4870 2884 4922
rect 2588 4868 2644 4870
rect 2668 4868 2724 4870
rect 2748 4868 2804 4870
rect 2828 4868 2884 4870
rect 2588 3834 2644 3836
rect 2668 3834 2724 3836
rect 2748 3834 2804 3836
rect 2828 3834 2884 3836
rect 2588 3782 2634 3834
rect 2634 3782 2644 3834
rect 2668 3782 2698 3834
rect 2698 3782 2710 3834
rect 2710 3782 2724 3834
rect 2748 3782 2762 3834
rect 2762 3782 2774 3834
rect 2774 3782 2804 3834
rect 2828 3782 2838 3834
rect 2838 3782 2884 3834
rect 2588 3780 2644 3782
rect 2668 3780 2724 3782
rect 2748 3780 2804 3782
rect 2828 3780 2884 3782
rect 7483 67482 7539 67484
rect 7563 67482 7619 67484
rect 7643 67482 7699 67484
rect 7723 67482 7779 67484
rect 7483 67430 7529 67482
rect 7529 67430 7539 67482
rect 7563 67430 7593 67482
rect 7593 67430 7605 67482
rect 7605 67430 7619 67482
rect 7643 67430 7657 67482
rect 7657 67430 7669 67482
rect 7669 67430 7699 67482
rect 7723 67430 7733 67482
rect 7733 67430 7779 67482
rect 7483 67428 7539 67430
rect 7563 67428 7619 67430
rect 7643 67428 7699 67430
rect 7723 67428 7779 67430
rect 7483 66394 7539 66396
rect 7563 66394 7619 66396
rect 7643 66394 7699 66396
rect 7723 66394 7779 66396
rect 7483 66342 7529 66394
rect 7529 66342 7539 66394
rect 7563 66342 7593 66394
rect 7593 66342 7605 66394
rect 7605 66342 7619 66394
rect 7643 66342 7657 66394
rect 7657 66342 7669 66394
rect 7669 66342 7699 66394
rect 7723 66342 7733 66394
rect 7733 66342 7779 66394
rect 7483 66340 7539 66342
rect 7563 66340 7619 66342
rect 7643 66340 7699 66342
rect 7723 66340 7779 66342
rect 7483 65306 7539 65308
rect 7563 65306 7619 65308
rect 7643 65306 7699 65308
rect 7723 65306 7779 65308
rect 7483 65254 7529 65306
rect 7529 65254 7539 65306
rect 7563 65254 7593 65306
rect 7593 65254 7605 65306
rect 7605 65254 7619 65306
rect 7643 65254 7657 65306
rect 7657 65254 7669 65306
rect 7669 65254 7699 65306
rect 7723 65254 7733 65306
rect 7733 65254 7779 65306
rect 7483 65252 7539 65254
rect 7563 65252 7619 65254
rect 7643 65252 7699 65254
rect 7723 65252 7779 65254
rect 7483 64218 7539 64220
rect 7563 64218 7619 64220
rect 7643 64218 7699 64220
rect 7723 64218 7779 64220
rect 7483 64166 7529 64218
rect 7529 64166 7539 64218
rect 7563 64166 7593 64218
rect 7593 64166 7605 64218
rect 7605 64166 7619 64218
rect 7643 64166 7657 64218
rect 7657 64166 7669 64218
rect 7669 64166 7699 64218
rect 7723 64166 7733 64218
rect 7733 64166 7779 64218
rect 7483 64164 7539 64166
rect 7563 64164 7619 64166
rect 7643 64164 7699 64166
rect 7723 64164 7779 64166
rect 7483 63130 7539 63132
rect 7563 63130 7619 63132
rect 7643 63130 7699 63132
rect 7723 63130 7779 63132
rect 7483 63078 7529 63130
rect 7529 63078 7539 63130
rect 7563 63078 7593 63130
rect 7593 63078 7605 63130
rect 7605 63078 7619 63130
rect 7643 63078 7657 63130
rect 7657 63078 7669 63130
rect 7669 63078 7699 63130
rect 7723 63078 7733 63130
rect 7733 63078 7779 63130
rect 7483 63076 7539 63078
rect 7563 63076 7619 63078
rect 7643 63076 7699 63078
rect 7723 63076 7779 63078
rect 7483 62042 7539 62044
rect 7563 62042 7619 62044
rect 7643 62042 7699 62044
rect 7723 62042 7779 62044
rect 7483 61990 7529 62042
rect 7529 61990 7539 62042
rect 7563 61990 7593 62042
rect 7593 61990 7605 62042
rect 7605 61990 7619 62042
rect 7643 61990 7657 62042
rect 7657 61990 7669 62042
rect 7669 61990 7699 62042
rect 7723 61990 7733 62042
rect 7733 61990 7779 62042
rect 7483 61988 7539 61990
rect 7563 61988 7619 61990
rect 7643 61988 7699 61990
rect 7723 61988 7779 61990
rect 7483 60954 7539 60956
rect 7563 60954 7619 60956
rect 7643 60954 7699 60956
rect 7723 60954 7779 60956
rect 7483 60902 7529 60954
rect 7529 60902 7539 60954
rect 7563 60902 7593 60954
rect 7593 60902 7605 60954
rect 7605 60902 7619 60954
rect 7643 60902 7657 60954
rect 7657 60902 7669 60954
rect 7669 60902 7699 60954
rect 7723 60902 7733 60954
rect 7733 60902 7779 60954
rect 7483 60900 7539 60902
rect 7563 60900 7619 60902
rect 7643 60900 7699 60902
rect 7723 60900 7779 60902
rect 7483 59866 7539 59868
rect 7563 59866 7619 59868
rect 7643 59866 7699 59868
rect 7723 59866 7779 59868
rect 7483 59814 7529 59866
rect 7529 59814 7539 59866
rect 7563 59814 7593 59866
rect 7593 59814 7605 59866
rect 7605 59814 7619 59866
rect 7643 59814 7657 59866
rect 7657 59814 7669 59866
rect 7669 59814 7699 59866
rect 7723 59814 7733 59866
rect 7733 59814 7779 59866
rect 7483 59812 7539 59814
rect 7563 59812 7619 59814
rect 7643 59812 7699 59814
rect 7723 59812 7779 59814
rect 7483 58778 7539 58780
rect 7563 58778 7619 58780
rect 7643 58778 7699 58780
rect 7723 58778 7779 58780
rect 7483 58726 7529 58778
rect 7529 58726 7539 58778
rect 7563 58726 7593 58778
rect 7593 58726 7605 58778
rect 7605 58726 7619 58778
rect 7643 58726 7657 58778
rect 7657 58726 7669 58778
rect 7669 58726 7699 58778
rect 7723 58726 7733 58778
rect 7733 58726 7779 58778
rect 7483 58724 7539 58726
rect 7563 58724 7619 58726
rect 7643 58724 7699 58726
rect 7723 58724 7779 58726
rect 7483 57690 7539 57692
rect 7563 57690 7619 57692
rect 7643 57690 7699 57692
rect 7723 57690 7779 57692
rect 7483 57638 7529 57690
rect 7529 57638 7539 57690
rect 7563 57638 7593 57690
rect 7593 57638 7605 57690
rect 7605 57638 7619 57690
rect 7643 57638 7657 57690
rect 7657 57638 7669 57690
rect 7669 57638 7699 57690
rect 7723 57638 7733 57690
rect 7733 57638 7779 57690
rect 7483 57636 7539 57638
rect 7563 57636 7619 57638
rect 7643 57636 7699 57638
rect 7723 57636 7779 57638
rect 7483 56602 7539 56604
rect 7563 56602 7619 56604
rect 7643 56602 7699 56604
rect 7723 56602 7779 56604
rect 7483 56550 7529 56602
rect 7529 56550 7539 56602
rect 7563 56550 7593 56602
rect 7593 56550 7605 56602
rect 7605 56550 7619 56602
rect 7643 56550 7657 56602
rect 7657 56550 7669 56602
rect 7669 56550 7699 56602
rect 7723 56550 7733 56602
rect 7733 56550 7779 56602
rect 7483 56548 7539 56550
rect 7563 56548 7619 56550
rect 7643 56548 7699 56550
rect 7723 56548 7779 56550
rect 7483 55514 7539 55516
rect 7563 55514 7619 55516
rect 7643 55514 7699 55516
rect 7723 55514 7779 55516
rect 7483 55462 7529 55514
rect 7529 55462 7539 55514
rect 7563 55462 7593 55514
rect 7593 55462 7605 55514
rect 7605 55462 7619 55514
rect 7643 55462 7657 55514
rect 7657 55462 7669 55514
rect 7669 55462 7699 55514
rect 7723 55462 7733 55514
rect 7733 55462 7779 55514
rect 7483 55460 7539 55462
rect 7563 55460 7619 55462
rect 7643 55460 7699 55462
rect 7723 55460 7779 55462
rect 7483 54426 7539 54428
rect 7563 54426 7619 54428
rect 7643 54426 7699 54428
rect 7723 54426 7779 54428
rect 7483 54374 7529 54426
rect 7529 54374 7539 54426
rect 7563 54374 7593 54426
rect 7593 54374 7605 54426
rect 7605 54374 7619 54426
rect 7643 54374 7657 54426
rect 7657 54374 7669 54426
rect 7669 54374 7699 54426
rect 7723 54374 7733 54426
rect 7733 54374 7779 54426
rect 7483 54372 7539 54374
rect 7563 54372 7619 54374
rect 7643 54372 7699 54374
rect 7723 54372 7779 54374
rect 7483 53338 7539 53340
rect 7563 53338 7619 53340
rect 7643 53338 7699 53340
rect 7723 53338 7779 53340
rect 7483 53286 7529 53338
rect 7529 53286 7539 53338
rect 7563 53286 7593 53338
rect 7593 53286 7605 53338
rect 7605 53286 7619 53338
rect 7643 53286 7657 53338
rect 7657 53286 7669 53338
rect 7669 53286 7699 53338
rect 7723 53286 7733 53338
rect 7733 53286 7779 53338
rect 7483 53284 7539 53286
rect 7563 53284 7619 53286
rect 7643 53284 7699 53286
rect 7723 53284 7779 53286
rect 7483 52250 7539 52252
rect 7563 52250 7619 52252
rect 7643 52250 7699 52252
rect 7723 52250 7779 52252
rect 7483 52198 7529 52250
rect 7529 52198 7539 52250
rect 7563 52198 7593 52250
rect 7593 52198 7605 52250
rect 7605 52198 7619 52250
rect 7643 52198 7657 52250
rect 7657 52198 7669 52250
rect 7669 52198 7699 52250
rect 7723 52198 7733 52250
rect 7733 52198 7779 52250
rect 7483 52196 7539 52198
rect 7563 52196 7619 52198
rect 7643 52196 7699 52198
rect 7723 52196 7779 52198
rect 7483 51162 7539 51164
rect 7563 51162 7619 51164
rect 7643 51162 7699 51164
rect 7723 51162 7779 51164
rect 7483 51110 7529 51162
rect 7529 51110 7539 51162
rect 7563 51110 7593 51162
rect 7593 51110 7605 51162
rect 7605 51110 7619 51162
rect 7643 51110 7657 51162
rect 7657 51110 7669 51162
rect 7669 51110 7699 51162
rect 7723 51110 7733 51162
rect 7733 51110 7779 51162
rect 7483 51108 7539 51110
rect 7563 51108 7619 51110
rect 7643 51108 7699 51110
rect 7723 51108 7779 51110
rect 7483 50074 7539 50076
rect 7563 50074 7619 50076
rect 7643 50074 7699 50076
rect 7723 50074 7779 50076
rect 7483 50022 7529 50074
rect 7529 50022 7539 50074
rect 7563 50022 7593 50074
rect 7593 50022 7605 50074
rect 7605 50022 7619 50074
rect 7643 50022 7657 50074
rect 7657 50022 7669 50074
rect 7669 50022 7699 50074
rect 7723 50022 7733 50074
rect 7733 50022 7779 50074
rect 7483 50020 7539 50022
rect 7563 50020 7619 50022
rect 7643 50020 7699 50022
rect 7723 50020 7779 50022
rect 7483 48986 7539 48988
rect 7563 48986 7619 48988
rect 7643 48986 7699 48988
rect 7723 48986 7779 48988
rect 7483 48934 7529 48986
rect 7529 48934 7539 48986
rect 7563 48934 7593 48986
rect 7593 48934 7605 48986
rect 7605 48934 7619 48986
rect 7643 48934 7657 48986
rect 7657 48934 7669 48986
rect 7669 48934 7699 48986
rect 7723 48934 7733 48986
rect 7733 48934 7779 48986
rect 7483 48932 7539 48934
rect 7563 48932 7619 48934
rect 7643 48932 7699 48934
rect 7723 48932 7779 48934
rect 7483 47898 7539 47900
rect 7563 47898 7619 47900
rect 7643 47898 7699 47900
rect 7723 47898 7779 47900
rect 7483 47846 7529 47898
rect 7529 47846 7539 47898
rect 7563 47846 7593 47898
rect 7593 47846 7605 47898
rect 7605 47846 7619 47898
rect 7643 47846 7657 47898
rect 7657 47846 7669 47898
rect 7669 47846 7699 47898
rect 7723 47846 7733 47898
rect 7733 47846 7779 47898
rect 7483 47844 7539 47846
rect 7563 47844 7619 47846
rect 7643 47844 7699 47846
rect 7723 47844 7779 47846
rect 7483 46810 7539 46812
rect 7563 46810 7619 46812
rect 7643 46810 7699 46812
rect 7723 46810 7779 46812
rect 7483 46758 7529 46810
rect 7529 46758 7539 46810
rect 7563 46758 7593 46810
rect 7593 46758 7605 46810
rect 7605 46758 7619 46810
rect 7643 46758 7657 46810
rect 7657 46758 7669 46810
rect 7669 46758 7699 46810
rect 7723 46758 7733 46810
rect 7733 46758 7779 46810
rect 7483 46756 7539 46758
rect 7563 46756 7619 46758
rect 7643 46756 7699 46758
rect 7723 46756 7779 46758
rect 7483 45722 7539 45724
rect 7563 45722 7619 45724
rect 7643 45722 7699 45724
rect 7723 45722 7779 45724
rect 7483 45670 7529 45722
rect 7529 45670 7539 45722
rect 7563 45670 7593 45722
rect 7593 45670 7605 45722
rect 7605 45670 7619 45722
rect 7643 45670 7657 45722
rect 7657 45670 7669 45722
rect 7669 45670 7699 45722
rect 7723 45670 7733 45722
rect 7733 45670 7779 45722
rect 7483 45668 7539 45670
rect 7563 45668 7619 45670
rect 7643 45668 7699 45670
rect 7723 45668 7779 45670
rect 7483 44634 7539 44636
rect 7563 44634 7619 44636
rect 7643 44634 7699 44636
rect 7723 44634 7779 44636
rect 7483 44582 7529 44634
rect 7529 44582 7539 44634
rect 7563 44582 7593 44634
rect 7593 44582 7605 44634
rect 7605 44582 7619 44634
rect 7643 44582 7657 44634
rect 7657 44582 7669 44634
rect 7669 44582 7699 44634
rect 7723 44582 7733 44634
rect 7733 44582 7779 44634
rect 7483 44580 7539 44582
rect 7563 44580 7619 44582
rect 7643 44580 7699 44582
rect 7723 44580 7779 44582
rect 7483 43546 7539 43548
rect 7563 43546 7619 43548
rect 7643 43546 7699 43548
rect 7723 43546 7779 43548
rect 7483 43494 7529 43546
rect 7529 43494 7539 43546
rect 7563 43494 7593 43546
rect 7593 43494 7605 43546
rect 7605 43494 7619 43546
rect 7643 43494 7657 43546
rect 7657 43494 7669 43546
rect 7669 43494 7699 43546
rect 7723 43494 7733 43546
rect 7733 43494 7779 43546
rect 7483 43492 7539 43494
rect 7563 43492 7619 43494
rect 7643 43492 7699 43494
rect 7723 43492 7779 43494
rect 7483 42458 7539 42460
rect 7563 42458 7619 42460
rect 7643 42458 7699 42460
rect 7723 42458 7779 42460
rect 7483 42406 7529 42458
rect 7529 42406 7539 42458
rect 7563 42406 7593 42458
rect 7593 42406 7605 42458
rect 7605 42406 7619 42458
rect 7643 42406 7657 42458
rect 7657 42406 7669 42458
rect 7669 42406 7699 42458
rect 7723 42406 7733 42458
rect 7733 42406 7779 42458
rect 7483 42404 7539 42406
rect 7563 42404 7619 42406
rect 7643 42404 7699 42406
rect 7723 42404 7779 42406
rect 7483 41370 7539 41372
rect 7563 41370 7619 41372
rect 7643 41370 7699 41372
rect 7723 41370 7779 41372
rect 7483 41318 7529 41370
rect 7529 41318 7539 41370
rect 7563 41318 7593 41370
rect 7593 41318 7605 41370
rect 7605 41318 7619 41370
rect 7643 41318 7657 41370
rect 7657 41318 7669 41370
rect 7669 41318 7699 41370
rect 7723 41318 7733 41370
rect 7733 41318 7779 41370
rect 7483 41316 7539 41318
rect 7563 41316 7619 41318
rect 7643 41316 7699 41318
rect 7723 41316 7779 41318
rect 7483 40282 7539 40284
rect 7563 40282 7619 40284
rect 7643 40282 7699 40284
rect 7723 40282 7779 40284
rect 7483 40230 7529 40282
rect 7529 40230 7539 40282
rect 7563 40230 7593 40282
rect 7593 40230 7605 40282
rect 7605 40230 7619 40282
rect 7643 40230 7657 40282
rect 7657 40230 7669 40282
rect 7669 40230 7699 40282
rect 7723 40230 7733 40282
rect 7733 40230 7779 40282
rect 7483 40228 7539 40230
rect 7563 40228 7619 40230
rect 7643 40228 7699 40230
rect 7723 40228 7779 40230
rect 7483 39194 7539 39196
rect 7563 39194 7619 39196
rect 7643 39194 7699 39196
rect 7723 39194 7779 39196
rect 7483 39142 7529 39194
rect 7529 39142 7539 39194
rect 7563 39142 7593 39194
rect 7593 39142 7605 39194
rect 7605 39142 7619 39194
rect 7643 39142 7657 39194
rect 7657 39142 7669 39194
rect 7669 39142 7699 39194
rect 7723 39142 7733 39194
rect 7733 39142 7779 39194
rect 7483 39140 7539 39142
rect 7563 39140 7619 39142
rect 7643 39140 7699 39142
rect 7723 39140 7779 39142
rect 7483 38106 7539 38108
rect 7563 38106 7619 38108
rect 7643 38106 7699 38108
rect 7723 38106 7779 38108
rect 7483 38054 7529 38106
rect 7529 38054 7539 38106
rect 7563 38054 7593 38106
rect 7593 38054 7605 38106
rect 7605 38054 7619 38106
rect 7643 38054 7657 38106
rect 7657 38054 7669 38106
rect 7669 38054 7699 38106
rect 7723 38054 7733 38106
rect 7733 38054 7779 38106
rect 7483 38052 7539 38054
rect 7563 38052 7619 38054
rect 7643 38052 7699 38054
rect 7723 38052 7779 38054
rect 7483 37018 7539 37020
rect 7563 37018 7619 37020
rect 7643 37018 7699 37020
rect 7723 37018 7779 37020
rect 7483 36966 7529 37018
rect 7529 36966 7539 37018
rect 7563 36966 7593 37018
rect 7593 36966 7605 37018
rect 7605 36966 7619 37018
rect 7643 36966 7657 37018
rect 7657 36966 7669 37018
rect 7669 36966 7699 37018
rect 7723 36966 7733 37018
rect 7733 36966 7779 37018
rect 7483 36964 7539 36966
rect 7563 36964 7619 36966
rect 7643 36964 7699 36966
rect 7723 36964 7779 36966
rect 7483 35930 7539 35932
rect 7563 35930 7619 35932
rect 7643 35930 7699 35932
rect 7723 35930 7779 35932
rect 7483 35878 7529 35930
rect 7529 35878 7539 35930
rect 7563 35878 7593 35930
rect 7593 35878 7605 35930
rect 7605 35878 7619 35930
rect 7643 35878 7657 35930
rect 7657 35878 7669 35930
rect 7669 35878 7699 35930
rect 7723 35878 7733 35930
rect 7733 35878 7779 35930
rect 7483 35876 7539 35878
rect 7563 35876 7619 35878
rect 7643 35876 7699 35878
rect 7723 35876 7779 35878
rect 7483 34842 7539 34844
rect 7563 34842 7619 34844
rect 7643 34842 7699 34844
rect 7723 34842 7779 34844
rect 7483 34790 7529 34842
rect 7529 34790 7539 34842
rect 7563 34790 7593 34842
rect 7593 34790 7605 34842
rect 7605 34790 7619 34842
rect 7643 34790 7657 34842
rect 7657 34790 7669 34842
rect 7669 34790 7699 34842
rect 7723 34790 7733 34842
rect 7733 34790 7779 34842
rect 7483 34788 7539 34790
rect 7563 34788 7619 34790
rect 7643 34788 7699 34790
rect 7723 34788 7779 34790
rect 7483 33754 7539 33756
rect 7563 33754 7619 33756
rect 7643 33754 7699 33756
rect 7723 33754 7779 33756
rect 7483 33702 7529 33754
rect 7529 33702 7539 33754
rect 7563 33702 7593 33754
rect 7593 33702 7605 33754
rect 7605 33702 7619 33754
rect 7643 33702 7657 33754
rect 7657 33702 7669 33754
rect 7669 33702 7699 33754
rect 7723 33702 7733 33754
rect 7733 33702 7779 33754
rect 7483 33700 7539 33702
rect 7563 33700 7619 33702
rect 7643 33700 7699 33702
rect 7723 33700 7779 33702
rect 7483 32666 7539 32668
rect 7563 32666 7619 32668
rect 7643 32666 7699 32668
rect 7723 32666 7779 32668
rect 7483 32614 7529 32666
rect 7529 32614 7539 32666
rect 7563 32614 7593 32666
rect 7593 32614 7605 32666
rect 7605 32614 7619 32666
rect 7643 32614 7657 32666
rect 7657 32614 7669 32666
rect 7669 32614 7699 32666
rect 7723 32614 7733 32666
rect 7733 32614 7779 32666
rect 7483 32612 7539 32614
rect 7563 32612 7619 32614
rect 7643 32612 7699 32614
rect 7723 32612 7779 32614
rect 7483 31578 7539 31580
rect 7563 31578 7619 31580
rect 7643 31578 7699 31580
rect 7723 31578 7779 31580
rect 7483 31526 7529 31578
rect 7529 31526 7539 31578
rect 7563 31526 7593 31578
rect 7593 31526 7605 31578
rect 7605 31526 7619 31578
rect 7643 31526 7657 31578
rect 7657 31526 7669 31578
rect 7669 31526 7699 31578
rect 7723 31526 7733 31578
rect 7733 31526 7779 31578
rect 7483 31524 7539 31526
rect 7563 31524 7619 31526
rect 7643 31524 7699 31526
rect 7723 31524 7779 31526
rect 7483 30490 7539 30492
rect 7563 30490 7619 30492
rect 7643 30490 7699 30492
rect 7723 30490 7779 30492
rect 7483 30438 7529 30490
rect 7529 30438 7539 30490
rect 7563 30438 7593 30490
rect 7593 30438 7605 30490
rect 7605 30438 7619 30490
rect 7643 30438 7657 30490
rect 7657 30438 7669 30490
rect 7669 30438 7699 30490
rect 7723 30438 7733 30490
rect 7733 30438 7779 30490
rect 7483 30436 7539 30438
rect 7563 30436 7619 30438
rect 7643 30436 7699 30438
rect 7723 30436 7779 30438
rect 7483 29402 7539 29404
rect 7563 29402 7619 29404
rect 7643 29402 7699 29404
rect 7723 29402 7779 29404
rect 7483 29350 7529 29402
rect 7529 29350 7539 29402
rect 7563 29350 7593 29402
rect 7593 29350 7605 29402
rect 7605 29350 7619 29402
rect 7643 29350 7657 29402
rect 7657 29350 7669 29402
rect 7669 29350 7699 29402
rect 7723 29350 7733 29402
rect 7733 29350 7779 29402
rect 7483 29348 7539 29350
rect 7563 29348 7619 29350
rect 7643 29348 7699 29350
rect 7723 29348 7779 29350
rect 7483 28314 7539 28316
rect 7563 28314 7619 28316
rect 7643 28314 7699 28316
rect 7723 28314 7779 28316
rect 7483 28262 7529 28314
rect 7529 28262 7539 28314
rect 7563 28262 7593 28314
rect 7593 28262 7605 28314
rect 7605 28262 7619 28314
rect 7643 28262 7657 28314
rect 7657 28262 7669 28314
rect 7669 28262 7699 28314
rect 7723 28262 7733 28314
rect 7733 28262 7779 28314
rect 7483 28260 7539 28262
rect 7563 28260 7619 28262
rect 7643 28260 7699 28262
rect 7723 28260 7779 28262
rect 7483 27226 7539 27228
rect 7563 27226 7619 27228
rect 7643 27226 7699 27228
rect 7723 27226 7779 27228
rect 7483 27174 7529 27226
rect 7529 27174 7539 27226
rect 7563 27174 7593 27226
rect 7593 27174 7605 27226
rect 7605 27174 7619 27226
rect 7643 27174 7657 27226
rect 7657 27174 7669 27226
rect 7669 27174 7699 27226
rect 7723 27174 7733 27226
rect 7733 27174 7779 27226
rect 7483 27172 7539 27174
rect 7563 27172 7619 27174
rect 7643 27172 7699 27174
rect 7723 27172 7779 27174
rect 7483 26138 7539 26140
rect 7563 26138 7619 26140
rect 7643 26138 7699 26140
rect 7723 26138 7779 26140
rect 7483 26086 7529 26138
rect 7529 26086 7539 26138
rect 7563 26086 7593 26138
rect 7593 26086 7605 26138
rect 7605 26086 7619 26138
rect 7643 26086 7657 26138
rect 7657 26086 7669 26138
rect 7669 26086 7699 26138
rect 7723 26086 7733 26138
rect 7733 26086 7779 26138
rect 7483 26084 7539 26086
rect 7563 26084 7619 26086
rect 7643 26084 7699 26086
rect 7723 26084 7779 26086
rect 7483 25050 7539 25052
rect 7563 25050 7619 25052
rect 7643 25050 7699 25052
rect 7723 25050 7779 25052
rect 7483 24998 7529 25050
rect 7529 24998 7539 25050
rect 7563 24998 7593 25050
rect 7593 24998 7605 25050
rect 7605 24998 7619 25050
rect 7643 24998 7657 25050
rect 7657 24998 7669 25050
rect 7669 24998 7699 25050
rect 7723 24998 7733 25050
rect 7733 24998 7779 25050
rect 7483 24996 7539 24998
rect 7563 24996 7619 24998
rect 7643 24996 7699 24998
rect 7723 24996 7779 24998
rect 7483 23962 7539 23964
rect 7563 23962 7619 23964
rect 7643 23962 7699 23964
rect 7723 23962 7779 23964
rect 7483 23910 7529 23962
rect 7529 23910 7539 23962
rect 7563 23910 7593 23962
rect 7593 23910 7605 23962
rect 7605 23910 7619 23962
rect 7643 23910 7657 23962
rect 7657 23910 7669 23962
rect 7669 23910 7699 23962
rect 7723 23910 7733 23962
rect 7733 23910 7779 23962
rect 7483 23908 7539 23910
rect 7563 23908 7619 23910
rect 7643 23908 7699 23910
rect 7723 23908 7779 23910
rect 7483 22874 7539 22876
rect 7563 22874 7619 22876
rect 7643 22874 7699 22876
rect 7723 22874 7779 22876
rect 7483 22822 7529 22874
rect 7529 22822 7539 22874
rect 7563 22822 7593 22874
rect 7593 22822 7605 22874
rect 7605 22822 7619 22874
rect 7643 22822 7657 22874
rect 7657 22822 7669 22874
rect 7669 22822 7699 22874
rect 7723 22822 7733 22874
rect 7733 22822 7779 22874
rect 7483 22820 7539 22822
rect 7563 22820 7619 22822
rect 7643 22820 7699 22822
rect 7723 22820 7779 22822
rect 7483 21786 7539 21788
rect 7563 21786 7619 21788
rect 7643 21786 7699 21788
rect 7723 21786 7779 21788
rect 7483 21734 7529 21786
rect 7529 21734 7539 21786
rect 7563 21734 7593 21786
rect 7593 21734 7605 21786
rect 7605 21734 7619 21786
rect 7643 21734 7657 21786
rect 7657 21734 7669 21786
rect 7669 21734 7699 21786
rect 7723 21734 7733 21786
rect 7733 21734 7779 21786
rect 7483 21732 7539 21734
rect 7563 21732 7619 21734
rect 7643 21732 7699 21734
rect 7723 21732 7779 21734
rect 7483 20698 7539 20700
rect 7563 20698 7619 20700
rect 7643 20698 7699 20700
rect 7723 20698 7779 20700
rect 7483 20646 7529 20698
rect 7529 20646 7539 20698
rect 7563 20646 7593 20698
rect 7593 20646 7605 20698
rect 7605 20646 7619 20698
rect 7643 20646 7657 20698
rect 7657 20646 7669 20698
rect 7669 20646 7699 20698
rect 7723 20646 7733 20698
rect 7733 20646 7779 20698
rect 7483 20644 7539 20646
rect 7563 20644 7619 20646
rect 7643 20644 7699 20646
rect 7723 20644 7779 20646
rect 7483 19610 7539 19612
rect 7563 19610 7619 19612
rect 7643 19610 7699 19612
rect 7723 19610 7779 19612
rect 7483 19558 7529 19610
rect 7529 19558 7539 19610
rect 7563 19558 7593 19610
rect 7593 19558 7605 19610
rect 7605 19558 7619 19610
rect 7643 19558 7657 19610
rect 7657 19558 7669 19610
rect 7669 19558 7699 19610
rect 7723 19558 7733 19610
rect 7733 19558 7779 19610
rect 7483 19556 7539 19558
rect 7563 19556 7619 19558
rect 7643 19556 7699 19558
rect 7723 19556 7779 19558
rect 10138 76064 10194 76120
rect 10138 74976 10194 75032
rect 9115 73466 9171 73468
rect 9195 73466 9251 73468
rect 9275 73466 9331 73468
rect 9355 73466 9411 73468
rect 9115 73414 9161 73466
rect 9161 73414 9171 73466
rect 9195 73414 9225 73466
rect 9225 73414 9237 73466
rect 9237 73414 9251 73466
rect 9275 73414 9289 73466
rect 9289 73414 9301 73466
rect 9301 73414 9331 73466
rect 9355 73414 9365 73466
rect 9365 73414 9411 73466
rect 9115 73412 9171 73414
rect 9195 73412 9251 73414
rect 9275 73412 9331 73414
rect 9355 73412 9411 73414
rect 10138 73888 10194 73944
rect 10138 72664 10194 72720
rect 9115 72378 9171 72380
rect 9195 72378 9251 72380
rect 9275 72378 9331 72380
rect 9355 72378 9411 72380
rect 9115 72326 9161 72378
rect 9161 72326 9171 72378
rect 9195 72326 9225 72378
rect 9225 72326 9237 72378
rect 9237 72326 9251 72378
rect 9275 72326 9289 72378
rect 9289 72326 9301 72378
rect 9301 72326 9331 72378
rect 9355 72326 9365 72378
rect 9365 72326 9411 72378
rect 9115 72324 9171 72326
rect 9195 72324 9251 72326
rect 9275 72324 9331 72326
rect 9355 72324 9411 72326
rect 10138 71576 10194 71632
rect 9115 71290 9171 71292
rect 9195 71290 9251 71292
rect 9275 71290 9331 71292
rect 9355 71290 9411 71292
rect 9115 71238 9161 71290
rect 9161 71238 9171 71290
rect 9195 71238 9225 71290
rect 9225 71238 9237 71290
rect 9237 71238 9251 71290
rect 9275 71238 9289 71290
rect 9289 71238 9301 71290
rect 9301 71238 9331 71290
rect 9355 71238 9365 71290
rect 9365 71238 9411 71290
rect 9115 71236 9171 71238
rect 9195 71236 9251 71238
rect 9275 71236 9331 71238
rect 9355 71236 9411 71238
rect 9115 70202 9171 70204
rect 9195 70202 9251 70204
rect 9275 70202 9331 70204
rect 9355 70202 9411 70204
rect 9115 70150 9161 70202
rect 9161 70150 9171 70202
rect 9195 70150 9225 70202
rect 9225 70150 9237 70202
rect 9237 70150 9251 70202
rect 9275 70150 9289 70202
rect 9289 70150 9301 70202
rect 9301 70150 9331 70202
rect 9355 70150 9365 70202
rect 9365 70150 9411 70202
rect 9115 70148 9171 70150
rect 9195 70148 9251 70150
rect 9275 70148 9331 70150
rect 9355 70148 9411 70150
rect 10138 70488 10194 70544
rect 10138 69400 10194 69456
rect 9115 69114 9171 69116
rect 9195 69114 9251 69116
rect 9275 69114 9331 69116
rect 9355 69114 9411 69116
rect 9115 69062 9161 69114
rect 9161 69062 9171 69114
rect 9195 69062 9225 69114
rect 9225 69062 9237 69114
rect 9237 69062 9251 69114
rect 9275 69062 9289 69114
rect 9289 69062 9301 69114
rect 9301 69062 9331 69114
rect 9355 69062 9365 69114
rect 9365 69062 9411 69114
rect 9115 69060 9171 69062
rect 9195 69060 9251 69062
rect 9275 69060 9331 69062
rect 9355 69060 9411 69062
rect 10138 68312 10194 68368
rect 9115 68026 9171 68028
rect 9195 68026 9251 68028
rect 9275 68026 9331 68028
rect 9355 68026 9411 68028
rect 9115 67974 9161 68026
rect 9161 67974 9171 68026
rect 9195 67974 9225 68026
rect 9225 67974 9237 68026
rect 9237 67974 9251 68026
rect 9275 67974 9289 68026
rect 9289 67974 9301 68026
rect 9301 67974 9331 68026
rect 9355 67974 9365 68026
rect 9365 67974 9411 68026
rect 9115 67972 9171 67974
rect 9195 67972 9251 67974
rect 9275 67972 9331 67974
rect 9355 67972 9411 67974
rect 9115 66938 9171 66940
rect 9195 66938 9251 66940
rect 9275 66938 9331 66940
rect 9355 66938 9411 66940
rect 9115 66886 9161 66938
rect 9161 66886 9171 66938
rect 9195 66886 9225 66938
rect 9225 66886 9237 66938
rect 9237 66886 9251 66938
rect 9275 66886 9289 66938
rect 9289 66886 9301 66938
rect 9301 66886 9331 66938
rect 9355 66886 9365 66938
rect 9365 66886 9411 66938
rect 9115 66884 9171 66886
rect 9195 66884 9251 66886
rect 9275 66884 9331 66886
rect 9355 66884 9411 66886
rect 10138 67224 10194 67280
rect 10138 66000 10194 66056
rect 9115 65850 9171 65852
rect 9195 65850 9251 65852
rect 9275 65850 9331 65852
rect 9355 65850 9411 65852
rect 9115 65798 9161 65850
rect 9161 65798 9171 65850
rect 9195 65798 9225 65850
rect 9225 65798 9237 65850
rect 9237 65798 9251 65850
rect 9275 65798 9289 65850
rect 9289 65798 9301 65850
rect 9301 65798 9331 65850
rect 9355 65798 9365 65850
rect 9365 65798 9411 65850
rect 9115 65796 9171 65798
rect 9195 65796 9251 65798
rect 9275 65796 9331 65798
rect 9355 65796 9411 65798
rect 10138 64912 10194 64968
rect 9115 64762 9171 64764
rect 9195 64762 9251 64764
rect 9275 64762 9331 64764
rect 9355 64762 9411 64764
rect 9115 64710 9161 64762
rect 9161 64710 9171 64762
rect 9195 64710 9225 64762
rect 9225 64710 9237 64762
rect 9237 64710 9251 64762
rect 9275 64710 9289 64762
rect 9289 64710 9301 64762
rect 9301 64710 9331 64762
rect 9355 64710 9365 64762
rect 9365 64710 9411 64762
rect 9115 64708 9171 64710
rect 9195 64708 9251 64710
rect 9275 64708 9331 64710
rect 9355 64708 9411 64710
rect 10138 63824 10194 63880
rect 9115 63674 9171 63676
rect 9195 63674 9251 63676
rect 9275 63674 9331 63676
rect 9355 63674 9411 63676
rect 9115 63622 9161 63674
rect 9161 63622 9171 63674
rect 9195 63622 9225 63674
rect 9225 63622 9237 63674
rect 9237 63622 9251 63674
rect 9275 63622 9289 63674
rect 9289 63622 9301 63674
rect 9301 63622 9331 63674
rect 9355 63622 9365 63674
rect 9365 63622 9411 63674
rect 9115 63620 9171 63622
rect 9195 63620 9251 63622
rect 9275 63620 9331 63622
rect 9355 63620 9411 63622
rect 10138 62736 10194 62792
rect 9115 62586 9171 62588
rect 9195 62586 9251 62588
rect 9275 62586 9331 62588
rect 9355 62586 9411 62588
rect 9115 62534 9161 62586
rect 9161 62534 9171 62586
rect 9195 62534 9225 62586
rect 9225 62534 9237 62586
rect 9237 62534 9251 62586
rect 9275 62534 9289 62586
rect 9289 62534 9301 62586
rect 9301 62534 9331 62586
rect 9355 62534 9365 62586
rect 9365 62534 9411 62586
rect 9115 62532 9171 62534
rect 9195 62532 9251 62534
rect 9275 62532 9331 62534
rect 9355 62532 9411 62534
rect 9115 61498 9171 61500
rect 9195 61498 9251 61500
rect 9275 61498 9331 61500
rect 9355 61498 9411 61500
rect 9115 61446 9161 61498
rect 9161 61446 9171 61498
rect 9195 61446 9225 61498
rect 9225 61446 9237 61498
rect 9237 61446 9251 61498
rect 9275 61446 9289 61498
rect 9289 61446 9301 61498
rect 9301 61446 9331 61498
rect 9355 61446 9365 61498
rect 9365 61446 9411 61498
rect 9115 61444 9171 61446
rect 9195 61444 9251 61446
rect 9275 61444 9331 61446
rect 9355 61444 9411 61446
rect 10138 61648 10194 61704
rect 10138 60560 10194 60616
rect 9115 60410 9171 60412
rect 9195 60410 9251 60412
rect 9275 60410 9331 60412
rect 9355 60410 9411 60412
rect 9115 60358 9161 60410
rect 9161 60358 9171 60410
rect 9195 60358 9225 60410
rect 9225 60358 9237 60410
rect 9237 60358 9251 60410
rect 9275 60358 9289 60410
rect 9289 60358 9301 60410
rect 9301 60358 9331 60410
rect 9355 60358 9365 60410
rect 9365 60358 9411 60410
rect 9115 60356 9171 60358
rect 9195 60356 9251 60358
rect 9275 60356 9331 60358
rect 9355 60356 9411 60358
rect 9115 59322 9171 59324
rect 9195 59322 9251 59324
rect 9275 59322 9331 59324
rect 9355 59322 9411 59324
rect 9115 59270 9161 59322
rect 9161 59270 9171 59322
rect 9195 59270 9225 59322
rect 9225 59270 9237 59322
rect 9237 59270 9251 59322
rect 9275 59270 9289 59322
rect 9289 59270 9301 59322
rect 9301 59270 9331 59322
rect 9355 59270 9365 59322
rect 9365 59270 9411 59322
rect 9115 59268 9171 59270
rect 9195 59268 9251 59270
rect 9275 59268 9331 59270
rect 9355 59268 9411 59270
rect 10138 59336 10194 59392
rect 10138 58248 10194 58304
rect 9115 58234 9171 58236
rect 9195 58234 9251 58236
rect 9275 58234 9331 58236
rect 9355 58234 9411 58236
rect 9115 58182 9161 58234
rect 9161 58182 9171 58234
rect 9195 58182 9225 58234
rect 9225 58182 9237 58234
rect 9237 58182 9251 58234
rect 9275 58182 9289 58234
rect 9289 58182 9301 58234
rect 9301 58182 9331 58234
rect 9355 58182 9365 58234
rect 9365 58182 9411 58234
rect 9115 58180 9171 58182
rect 9195 58180 9251 58182
rect 9275 58180 9331 58182
rect 9355 58180 9411 58182
rect 9115 57146 9171 57148
rect 9195 57146 9251 57148
rect 9275 57146 9331 57148
rect 9355 57146 9411 57148
rect 9115 57094 9161 57146
rect 9161 57094 9171 57146
rect 9195 57094 9225 57146
rect 9225 57094 9237 57146
rect 9237 57094 9251 57146
rect 9275 57094 9289 57146
rect 9289 57094 9301 57146
rect 9301 57094 9331 57146
rect 9355 57094 9365 57146
rect 9365 57094 9411 57146
rect 9115 57092 9171 57094
rect 9195 57092 9251 57094
rect 9275 57092 9331 57094
rect 9355 57092 9411 57094
rect 9115 56058 9171 56060
rect 9195 56058 9251 56060
rect 9275 56058 9331 56060
rect 9355 56058 9411 56060
rect 9115 56006 9161 56058
rect 9161 56006 9171 56058
rect 9195 56006 9225 56058
rect 9225 56006 9237 56058
rect 9237 56006 9251 56058
rect 9275 56006 9289 56058
rect 9289 56006 9301 56058
rect 9301 56006 9331 56058
rect 9355 56006 9365 56058
rect 9365 56006 9411 56058
rect 9115 56004 9171 56006
rect 9195 56004 9251 56006
rect 9275 56004 9331 56006
rect 9355 56004 9411 56006
rect 10138 57160 10194 57216
rect 10138 56072 10194 56128
rect 10138 54984 10194 55040
rect 9115 54970 9171 54972
rect 9195 54970 9251 54972
rect 9275 54970 9331 54972
rect 9355 54970 9411 54972
rect 9115 54918 9161 54970
rect 9161 54918 9171 54970
rect 9195 54918 9225 54970
rect 9225 54918 9237 54970
rect 9237 54918 9251 54970
rect 9275 54918 9289 54970
rect 9289 54918 9301 54970
rect 9301 54918 9331 54970
rect 9355 54918 9365 54970
rect 9365 54918 9411 54970
rect 9115 54916 9171 54918
rect 9195 54916 9251 54918
rect 9275 54916 9331 54918
rect 9355 54916 9411 54918
rect 9115 53882 9171 53884
rect 9195 53882 9251 53884
rect 9275 53882 9331 53884
rect 9355 53882 9411 53884
rect 9115 53830 9161 53882
rect 9161 53830 9171 53882
rect 9195 53830 9225 53882
rect 9225 53830 9237 53882
rect 9237 53830 9251 53882
rect 9275 53830 9289 53882
rect 9289 53830 9301 53882
rect 9301 53830 9331 53882
rect 9355 53830 9365 53882
rect 9365 53830 9411 53882
rect 9115 53828 9171 53830
rect 9195 53828 9251 53830
rect 9275 53828 9331 53830
rect 9355 53828 9411 53830
rect 10138 53896 10194 53952
rect 9115 52794 9171 52796
rect 9195 52794 9251 52796
rect 9275 52794 9331 52796
rect 9355 52794 9411 52796
rect 9115 52742 9161 52794
rect 9161 52742 9171 52794
rect 9195 52742 9225 52794
rect 9225 52742 9237 52794
rect 9237 52742 9251 52794
rect 9275 52742 9289 52794
rect 9289 52742 9301 52794
rect 9301 52742 9331 52794
rect 9355 52742 9365 52794
rect 9365 52742 9411 52794
rect 9115 52740 9171 52742
rect 9195 52740 9251 52742
rect 9275 52740 9331 52742
rect 9355 52740 9411 52742
rect 10138 52672 10194 52728
rect 9115 51706 9171 51708
rect 9195 51706 9251 51708
rect 9275 51706 9331 51708
rect 9355 51706 9411 51708
rect 9115 51654 9161 51706
rect 9161 51654 9171 51706
rect 9195 51654 9225 51706
rect 9225 51654 9237 51706
rect 9237 51654 9251 51706
rect 9275 51654 9289 51706
rect 9289 51654 9301 51706
rect 9301 51654 9331 51706
rect 9355 51654 9365 51706
rect 9365 51654 9411 51706
rect 9115 51652 9171 51654
rect 9195 51652 9251 51654
rect 9275 51652 9331 51654
rect 9355 51652 9411 51654
rect 10138 51584 10194 51640
rect 9115 50618 9171 50620
rect 9195 50618 9251 50620
rect 9275 50618 9331 50620
rect 9355 50618 9411 50620
rect 9115 50566 9161 50618
rect 9161 50566 9171 50618
rect 9195 50566 9225 50618
rect 9225 50566 9237 50618
rect 9237 50566 9251 50618
rect 9275 50566 9289 50618
rect 9289 50566 9301 50618
rect 9301 50566 9331 50618
rect 9355 50566 9365 50618
rect 9365 50566 9411 50618
rect 9115 50564 9171 50566
rect 9195 50564 9251 50566
rect 9275 50564 9331 50566
rect 9355 50564 9411 50566
rect 10138 50496 10194 50552
rect 9115 49530 9171 49532
rect 9195 49530 9251 49532
rect 9275 49530 9331 49532
rect 9355 49530 9411 49532
rect 9115 49478 9161 49530
rect 9161 49478 9171 49530
rect 9195 49478 9225 49530
rect 9225 49478 9237 49530
rect 9237 49478 9251 49530
rect 9275 49478 9289 49530
rect 9289 49478 9301 49530
rect 9301 49478 9331 49530
rect 9355 49478 9365 49530
rect 9365 49478 9411 49530
rect 9115 49476 9171 49478
rect 9195 49476 9251 49478
rect 9275 49476 9331 49478
rect 9355 49476 9411 49478
rect 10138 49408 10194 49464
rect 9115 48442 9171 48444
rect 9195 48442 9251 48444
rect 9275 48442 9331 48444
rect 9355 48442 9411 48444
rect 9115 48390 9161 48442
rect 9161 48390 9171 48442
rect 9195 48390 9225 48442
rect 9225 48390 9237 48442
rect 9237 48390 9251 48442
rect 9275 48390 9289 48442
rect 9289 48390 9301 48442
rect 9301 48390 9331 48442
rect 9355 48390 9365 48442
rect 9365 48390 9411 48442
rect 9115 48388 9171 48390
rect 9195 48388 9251 48390
rect 9275 48388 9331 48390
rect 9355 48388 9411 48390
rect 10138 48320 10194 48376
rect 9115 47354 9171 47356
rect 9195 47354 9251 47356
rect 9275 47354 9331 47356
rect 9355 47354 9411 47356
rect 9115 47302 9161 47354
rect 9161 47302 9171 47354
rect 9195 47302 9225 47354
rect 9225 47302 9237 47354
rect 9237 47302 9251 47354
rect 9275 47302 9289 47354
rect 9289 47302 9301 47354
rect 9301 47302 9331 47354
rect 9355 47302 9365 47354
rect 9365 47302 9411 47354
rect 9115 47300 9171 47302
rect 9195 47300 9251 47302
rect 9275 47300 9331 47302
rect 9355 47300 9411 47302
rect 10138 47232 10194 47288
rect 9115 46266 9171 46268
rect 9195 46266 9251 46268
rect 9275 46266 9331 46268
rect 9355 46266 9411 46268
rect 9115 46214 9161 46266
rect 9161 46214 9171 46266
rect 9195 46214 9225 46266
rect 9225 46214 9237 46266
rect 9237 46214 9251 46266
rect 9275 46214 9289 46266
rect 9289 46214 9301 46266
rect 9301 46214 9331 46266
rect 9355 46214 9365 46266
rect 9365 46214 9411 46266
rect 9115 46212 9171 46214
rect 9195 46212 9251 46214
rect 9275 46212 9331 46214
rect 9355 46212 9411 46214
rect 9115 45178 9171 45180
rect 9195 45178 9251 45180
rect 9275 45178 9331 45180
rect 9355 45178 9411 45180
rect 9115 45126 9161 45178
rect 9161 45126 9171 45178
rect 9195 45126 9225 45178
rect 9225 45126 9237 45178
rect 9237 45126 9251 45178
rect 9275 45126 9289 45178
rect 9289 45126 9301 45178
rect 9301 45126 9331 45178
rect 9355 45126 9365 45178
rect 9365 45126 9411 45178
rect 9115 45124 9171 45126
rect 9195 45124 9251 45126
rect 9275 45124 9331 45126
rect 9355 45124 9411 45126
rect 9115 44090 9171 44092
rect 9195 44090 9251 44092
rect 9275 44090 9331 44092
rect 9355 44090 9411 44092
rect 9115 44038 9161 44090
rect 9161 44038 9171 44090
rect 9195 44038 9225 44090
rect 9225 44038 9237 44090
rect 9237 44038 9251 44090
rect 9275 44038 9289 44090
rect 9289 44038 9301 44090
rect 9301 44038 9331 44090
rect 9355 44038 9365 44090
rect 9365 44038 9411 44090
rect 9115 44036 9171 44038
rect 9195 44036 9251 44038
rect 9275 44036 9331 44038
rect 9355 44036 9411 44038
rect 10138 46008 10194 46064
rect 10138 44920 10194 44976
rect 10138 43832 10194 43888
rect 9115 43002 9171 43004
rect 9195 43002 9251 43004
rect 9275 43002 9331 43004
rect 9355 43002 9411 43004
rect 9115 42950 9161 43002
rect 9161 42950 9171 43002
rect 9195 42950 9225 43002
rect 9225 42950 9237 43002
rect 9237 42950 9251 43002
rect 9275 42950 9289 43002
rect 9289 42950 9301 43002
rect 9301 42950 9331 43002
rect 9355 42950 9365 43002
rect 9365 42950 9411 43002
rect 9115 42948 9171 42950
rect 9195 42948 9251 42950
rect 9275 42948 9331 42950
rect 9355 42948 9411 42950
rect 10046 42744 10102 42800
rect 9115 41914 9171 41916
rect 9195 41914 9251 41916
rect 9275 41914 9331 41916
rect 9355 41914 9411 41916
rect 9115 41862 9161 41914
rect 9161 41862 9171 41914
rect 9195 41862 9225 41914
rect 9225 41862 9237 41914
rect 9237 41862 9251 41914
rect 9275 41862 9289 41914
rect 9289 41862 9301 41914
rect 9301 41862 9331 41914
rect 9355 41862 9365 41914
rect 9365 41862 9411 41914
rect 9115 41860 9171 41862
rect 9195 41860 9251 41862
rect 9275 41860 9331 41862
rect 9355 41860 9411 41862
rect 10046 41656 10102 41712
rect 9115 40826 9171 40828
rect 9195 40826 9251 40828
rect 9275 40826 9331 40828
rect 9355 40826 9411 40828
rect 9115 40774 9161 40826
rect 9161 40774 9171 40826
rect 9195 40774 9225 40826
rect 9225 40774 9237 40826
rect 9237 40774 9251 40826
rect 9275 40774 9289 40826
rect 9289 40774 9301 40826
rect 9301 40774 9331 40826
rect 9355 40774 9365 40826
rect 9365 40774 9411 40826
rect 9115 40772 9171 40774
rect 9195 40772 9251 40774
rect 9275 40772 9331 40774
rect 9355 40772 9411 40774
rect 10046 40568 10102 40624
rect 9115 39738 9171 39740
rect 9195 39738 9251 39740
rect 9275 39738 9331 39740
rect 9355 39738 9411 39740
rect 9115 39686 9161 39738
rect 9161 39686 9171 39738
rect 9195 39686 9225 39738
rect 9225 39686 9237 39738
rect 9237 39686 9251 39738
rect 9275 39686 9289 39738
rect 9289 39686 9301 39738
rect 9301 39686 9331 39738
rect 9355 39686 9365 39738
rect 9365 39686 9411 39738
rect 9115 39684 9171 39686
rect 9195 39684 9251 39686
rect 9275 39684 9331 39686
rect 9355 39684 9411 39686
rect 10046 39344 10102 39400
rect 9115 38650 9171 38652
rect 9195 38650 9251 38652
rect 9275 38650 9331 38652
rect 9355 38650 9411 38652
rect 9115 38598 9161 38650
rect 9161 38598 9171 38650
rect 9195 38598 9225 38650
rect 9225 38598 9237 38650
rect 9237 38598 9251 38650
rect 9275 38598 9289 38650
rect 9289 38598 9301 38650
rect 9301 38598 9331 38650
rect 9355 38598 9365 38650
rect 9365 38598 9411 38650
rect 9115 38596 9171 38598
rect 9195 38596 9251 38598
rect 9275 38596 9331 38598
rect 9355 38596 9411 38598
rect 10046 38256 10102 38312
rect 9115 37562 9171 37564
rect 9195 37562 9251 37564
rect 9275 37562 9331 37564
rect 9355 37562 9411 37564
rect 9115 37510 9161 37562
rect 9161 37510 9171 37562
rect 9195 37510 9225 37562
rect 9225 37510 9237 37562
rect 9237 37510 9251 37562
rect 9275 37510 9289 37562
rect 9289 37510 9301 37562
rect 9301 37510 9331 37562
rect 9355 37510 9365 37562
rect 9365 37510 9411 37562
rect 9115 37508 9171 37510
rect 9195 37508 9251 37510
rect 9275 37508 9331 37510
rect 9355 37508 9411 37510
rect 10046 37168 10102 37224
rect 9115 36474 9171 36476
rect 9195 36474 9251 36476
rect 9275 36474 9331 36476
rect 9355 36474 9411 36476
rect 9115 36422 9161 36474
rect 9161 36422 9171 36474
rect 9195 36422 9225 36474
rect 9225 36422 9237 36474
rect 9237 36422 9251 36474
rect 9275 36422 9289 36474
rect 9289 36422 9301 36474
rect 9301 36422 9331 36474
rect 9355 36422 9365 36474
rect 9365 36422 9411 36474
rect 9115 36420 9171 36422
rect 9195 36420 9251 36422
rect 9275 36420 9331 36422
rect 9355 36420 9411 36422
rect 10046 36080 10102 36136
rect 9115 35386 9171 35388
rect 9195 35386 9251 35388
rect 9275 35386 9331 35388
rect 9355 35386 9411 35388
rect 9115 35334 9161 35386
rect 9161 35334 9171 35386
rect 9195 35334 9225 35386
rect 9225 35334 9237 35386
rect 9237 35334 9251 35386
rect 9275 35334 9289 35386
rect 9289 35334 9301 35386
rect 9301 35334 9331 35386
rect 9355 35334 9365 35386
rect 9365 35334 9411 35386
rect 9115 35332 9171 35334
rect 9195 35332 9251 35334
rect 9275 35332 9331 35334
rect 9355 35332 9411 35334
rect 10046 34992 10102 35048
rect 9115 34298 9171 34300
rect 9195 34298 9251 34300
rect 9275 34298 9331 34300
rect 9355 34298 9411 34300
rect 9115 34246 9161 34298
rect 9161 34246 9171 34298
rect 9195 34246 9225 34298
rect 9225 34246 9237 34298
rect 9237 34246 9251 34298
rect 9275 34246 9289 34298
rect 9289 34246 9301 34298
rect 9301 34246 9331 34298
rect 9355 34246 9365 34298
rect 9365 34246 9411 34298
rect 9115 34244 9171 34246
rect 9195 34244 9251 34246
rect 9275 34244 9331 34246
rect 9355 34244 9411 34246
rect 10046 33904 10102 33960
rect 9115 33210 9171 33212
rect 9195 33210 9251 33212
rect 9275 33210 9331 33212
rect 9355 33210 9411 33212
rect 9115 33158 9161 33210
rect 9161 33158 9171 33210
rect 9195 33158 9225 33210
rect 9225 33158 9237 33210
rect 9237 33158 9251 33210
rect 9275 33158 9289 33210
rect 9289 33158 9301 33210
rect 9301 33158 9331 33210
rect 9355 33158 9365 33210
rect 9365 33158 9411 33210
rect 9115 33156 9171 33158
rect 9195 33156 9251 33158
rect 9275 33156 9331 33158
rect 9355 33156 9411 33158
rect 10046 32716 10048 32736
rect 10048 32716 10100 32736
rect 10100 32716 10102 32736
rect 10046 32680 10102 32716
rect 9115 32122 9171 32124
rect 9195 32122 9251 32124
rect 9275 32122 9331 32124
rect 9355 32122 9411 32124
rect 9115 32070 9161 32122
rect 9161 32070 9171 32122
rect 9195 32070 9225 32122
rect 9225 32070 9237 32122
rect 9237 32070 9251 32122
rect 9275 32070 9289 32122
rect 9289 32070 9301 32122
rect 9301 32070 9331 32122
rect 9355 32070 9365 32122
rect 9365 32070 9411 32122
rect 9115 32068 9171 32070
rect 9195 32068 9251 32070
rect 9275 32068 9331 32070
rect 9355 32068 9411 32070
rect 10046 31628 10048 31648
rect 10048 31628 10100 31648
rect 10100 31628 10102 31648
rect 10046 31592 10102 31628
rect 9115 31034 9171 31036
rect 9195 31034 9251 31036
rect 9275 31034 9331 31036
rect 9355 31034 9411 31036
rect 9115 30982 9161 31034
rect 9161 30982 9171 31034
rect 9195 30982 9225 31034
rect 9225 30982 9237 31034
rect 9237 30982 9251 31034
rect 9275 30982 9289 31034
rect 9289 30982 9301 31034
rect 9301 30982 9331 31034
rect 9355 30982 9365 31034
rect 9365 30982 9411 31034
rect 9115 30980 9171 30982
rect 9195 30980 9251 30982
rect 9275 30980 9331 30982
rect 9355 30980 9411 30982
rect 10046 30540 10048 30560
rect 10048 30540 10100 30560
rect 10100 30540 10102 30560
rect 9115 29946 9171 29948
rect 9195 29946 9251 29948
rect 9275 29946 9331 29948
rect 9355 29946 9411 29948
rect 9115 29894 9161 29946
rect 9161 29894 9171 29946
rect 9195 29894 9225 29946
rect 9225 29894 9237 29946
rect 9237 29894 9251 29946
rect 9275 29894 9289 29946
rect 9289 29894 9301 29946
rect 9301 29894 9331 29946
rect 9355 29894 9365 29946
rect 9365 29894 9411 29946
rect 9115 29892 9171 29894
rect 9195 29892 9251 29894
rect 9275 29892 9331 29894
rect 9355 29892 9411 29894
rect 10046 30504 10102 30540
rect 10046 29452 10048 29472
rect 10048 29452 10100 29472
rect 10100 29452 10102 29472
rect 10046 29416 10102 29452
rect 9115 28858 9171 28860
rect 9195 28858 9251 28860
rect 9275 28858 9331 28860
rect 9355 28858 9411 28860
rect 9115 28806 9161 28858
rect 9161 28806 9171 28858
rect 9195 28806 9225 28858
rect 9225 28806 9237 28858
rect 9237 28806 9251 28858
rect 9275 28806 9289 28858
rect 9289 28806 9301 28858
rect 9301 28806 9331 28858
rect 9355 28806 9365 28858
rect 9365 28806 9411 28858
rect 9115 28804 9171 28806
rect 9195 28804 9251 28806
rect 9275 28804 9331 28806
rect 9355 28804 9411 28806
rect 10046 28364 10048 28384
rect 10048 28364 10100 28384
rect 10100 28364 10102 28384
rect 10046 28328 10102 28364
rect 9115 27770 9171 27772
rect 9195 27770 9251 27772
rect 9275 27770 9331 27772
rect 9355 27770 9411 27772
rect 9115 27718 9161 27770
rect 9161 27718 9171 27770
rect 9195 27718 9225 27770
rect 9225 27718 9237 27770
rect 9237 27718 9251 27770
rect 9275 27718 9289 27770
rect 9289 27718 9301 27770
rect 9301 27718 9331 27770
rect 9355 27718 9365 27770
rect 9365 27718 9411 27770
rect 9115 27716 9171 27718
rect 9195 27716 9251 27718
rect 9275 27716 9331 27718
rect 9355 27716 9411 27718
rect 10046 27276 10048 27296
rect 10048 27276 10100 27296
rect 10100 27276 10102 27296
rect 10046 27240 10102 27276
rect 9115 26682 9171 26684
rect 9195 26682 9251 26684
rect 9275 26682 9331 26684
rect 9355 26682 9411 26684
rect 9115 26630 9161 26682
rect 9161 26630 9171 26682
rect 9195 26630 9225 26682
rect 9225 26630 9237 26682
rect 9237 26630 9251 26682
rect 9275 26630 9289 26682
rect 9289 26630 9301 26682
rect 9301 26630 9331 26682
rect 9355 26630 9365 26682
rect 9365 26630 9411 26682
rect 9115 26628 9171 26630
rect 9195 26628 9251 26630
rect 9275 26628 9331 26630
rect 9355 26628 9411 26630
rect 9115 25594 9171 25596
rect 9195 25594 9251 25596
rect 9275 25594 9331 25596
rect 9355 25594 9411 25596
rect 9115 25542 9161 25594
rect 9161 25542 9171 25594
rect 9195 25542 9225 25594
rect 9225 25542 9237 25594
rect 9237 25542 9251 25594
rect 9275 25542 9289 25594
rect 9289 25542 9301 25594
rect 9301 25542 9331 25594
rect 9355 25542 9365 25594
rect 9365 25542 9411 25594
rect 9115 25540 9171 25542
rect 9195 25540 9251 25542
rect 9275 25540 9331 25542
rect 9355 25540 9411 25542
rect 9115 24506 9171 24508
rect 9195 24506 9251 24508
rect 9275 24506 9331 24508
rect 9355 24506 9411 24508
rect 9115 24454 9161 24506
rect 9161 24454 9171 24506
rect 9195 24454 9225 24506
rect 9225 24454 9237 24506
rect 9237 24454 9251 24506
rect 9275 24454 9289 24506
rect 9289 24454 9301 24506
rect 9301 24454 9331 24506
rect 9355 24454 9365 24506
rect 9365 24454 9411 24506
rect 9115 24452 9171 24454
rect 9195 24452 9251 24454
rect 9275 24452 9331 24454
rect 9355 24452 9411 24454
rect 10046 26016 10102 26072
rect 10046 24928 10102 24984
rect 10046 23840 10102 23896
rect 9115 23418 9171 23420
rect 9195 23418 9251 23420
rect 9275 23418 9331 23420
rect 9355 23418 9411 23420
rect 9115 23366 9161 23418
rect 9161 23366 9171 23418
rect 9195 23366 9225 23418
rect 9225 23366 9237 23418
rect 9237 23366 9251 23418
rect 9275 23366 9289 23418
rect 9289 23366 9301 23418
rect 9301 23366 9331 23418
rect 9355 23366 9365 23418
rect 9365 23366 9411 23418
rect 9115 23364 9171 23366
rect 9195 23364 9251 23366
rect 9275 23364 9331 23366
rect 9355 23364 9411 23366
rect 10046 22752 10102 22808
rect 9115 22330 9171 22332
rect 9195 22330 9251 22332
rect 9275 22330 9331 22332
rect 9355 22330 9411 22332
rect 9115 22278 9161 22330
rect 9161 22278 9171 22330
rect 9195 22278 9225 22330
rect 9225 22278 9237 22330
rect 9237 22278 9251 22330
rect 9275 22278 9289 22330
rect 9289 22278 9301 22330
rect 9301 22278 9331 22330
rect 9355 22278 9365 22330
rect 9365 22278 9411 22330
rect 9115 22276 9171 22278
rect 9195 22276 9251 22278
rect 9275 22276 9331 22278
rect 9355 22276 9411 22278
rect 9115 21242 9171 21244
rect 9195 21242 9251 21244
rect 9275 21242 9331 21244
rect 9355 21242 9411 21244
rect 9115 21190 9161 21242
rect 9161 21190 9171 21242
rect 9195 21190 9225 21242
rect 9225 21190 9237 21242
rect 9237 21190 9251 21242
rect 9275 21190 9289 21242
rect 9289 21190 9301 21242
rect 9301 21190 9331 21242
rect 9355 21190 9365 21242
rect 9365 21190 9411 21242
rect 9115 21188 9171 21190
rect 9195 21188 9251 21190
rect 9275 21188 9331 21190
rect 9355 21188 9411 21190
rect 9115 20154 9171 20156
rect 9195 20154 9251 20156
rect 9275 20154 9331 20156
rect 9355 20154 9411 20156
rect 9115 20102 9161 20154
rect 9161 20102 9171 20154
rect 9195 20102 9225 20154
rect 9225 20102 9237 20154
rect 9237 20102 9251 20154
rect 9275 20102 9289 20154
rect 9289 20102 9301 20154
rect 9301 20102 9331 20154
rect 9355 20102 9365 20154
rect 9365 20102 9411 20154
rect 9115 20100 9171 20102
rect 9195 20100 9251 20102
rect 9275 20100 9331 20102
rect 9355 20100 9411 20102
rect 10046 21664 10102 21720
rect 10046 20576 10102 20632
rect 10046 19352 10102 19408
rect 9115 19066 9171 19068
rect 9195 19066 9251 19068
rect 9275 19066 9331 19068
rect 9355 19066 9411 19068
rect 9115 19014 9161 19066
rect 9161 19014 9171 19066
rect 9195 19014 9225 19066
rect 9225 19014 9237 19066
rect 9237 19014 9251 19066
rect 9275 19014 9289 19066
rect 9289 19014 9301 19066
rect 9301 19014 9331 19066
rect 9355 19014 9365 19066
rect 9365 19014 9411 19066
rect 9115 19012 9171 19014
rect 9195 19012 9251 19014
rect 9275 19012 9331 19014
rect 9355 19012 9411 19014
rect 7483 18522 7539 18524
rect 7563 18522 7619 18524
rect 7643 18522 7699 18524
rect 7723 18522 7779 18524
rect 7483 18470 7529 18522
rect 7529 18470 7539 18522
rect 7563 18470 7593 18522
rect 7593 18470 7605 18522
rect 7605 18470 7619 18522
rect 7643 18470 7657 18522
rect 7657 18470 7669 18522
rect 7669 18470 7699 18522
rect 7723 18470 7733 18522
rect 7733 18470 7779 18522
rect 7483 18468 7539 18470
rect 7563 18468 7619 18470
rect 7643 18468 7699 18470
rect 7723 18468 7779 18470
rect 10046 18264 10102 18320
rect 9115 17978 9171 17980
rect 9195 17978 9251 17980
rect 9275 17978 9331 17980
rect 9355 17978 9411 17980
rect 9115 17926 9161 17978
rect 9161 17926 9171 17978
rect 9195 17926 9225 17978
rect 9225 17926 9237 17978
rect 9237 17926 9251 17978
rect 9275 17926 9289 17978
rect 9289 17926 9301 17978
rect 9301 17926 9331 17978
rect 9355 17926 9365 17978
rect 9365 17926 9411 17978
rect 9115 17924 9171 17926
rect 9195 17924 9251 17926
rect 9275 17924 9331 17926
rect 9355 17924 9411 17926
rect 7483 17434 7539 17436
rect 7563 17434 7619 17436
rect 7643 17434 7699 17436
rect 7723 17434 7779 17436
rect 7483 17382 7529 17434
rect 7529 17382 7539 17434
rect 7563 17382 7593 17434
rect 7593 17382 7605 17434
rect 7605 17382 7619 17434
rect 7643 17382 7657 17434
rect 7657 17382 7669 17434
rect 7669 17382 7699 17434
rect 7723 17382 7733 17434
rect 7733 17382 7779 17434
rect 7483 17380 7539 17382
rect 7563 17380 7619 17382
rect 7643 17380 7699 17382
rect 7723 17380 7779 17382
rect 9115 16890 9171 16892
rect 9195 16890 9251 16892
rect 9275 16890 9331 16892
rect 9355 16890 9411 16892
rect 9115 16838 9161 16890
rect 9161 16838 9171 16890
rect 9195 16838 9225 16890
rect 9225 16838 9237 16890
rect 9237 16838 9251 16890
rect 9275 16838 9289 16890
rect 9289 16838 9301 16890
rect 9301 16838 9331 16890
rect 9355 16838 9365 16890
rect 9365 16838 9411 16890
rect 9115 16836 9171 16838
rect 9195 16836 9251 16838
rect 9275 16836 9331 16838
rect 9355 16836 9411 16838
rect 10046 17176 10102 17232
rect 7483 16346 7539 16348
rect 7563 16346 7619 16348
rect 7643 16346 7699 16348
rect 7723 16346 7779 16348
rect 7483 16294 7529 16346
rect 7529 16294 7539 16346
rect 7563 16294 7593 16346
rect 7593 16294 7605 16346
rect 7605 16294 7619 16346
rect 7643 16294 7657 16346
rect 7657 16294 7669 16346
rect 7669 16294 7699 16346
rect 7723 16294 7733 16346
rect 7733 16294 7779 16346
rect 7483 16292 7539 16294
rect 7563 16292 7619 16294
rect 7643 16292 7699 16294
rect 7723 16292 7779 16294
rect 9115 15802 9171 15804
rect 9195 15802 9251 15804
rect 9275 15802 9331 15804
rect 9355 15802 9411 15804
rect 9115 15750 9161 15802
rect 9161 15750 9171 15802
rect 9195 15750 9225 15802
rect 9225 15750 9237 15802
rect 9237 15750 9251 15802
rect 9275 15750 9289 15802
rect 9289 15750 9301 15802
rect 9301 15750 9331 15802
rect 9355 15750 9365 15802
rect 9365 15750 9411 15802
rect 9115 15748 9171 15750
rect 9195 15748 9251 15750
rect 9275 15748 9331 15750
rect 9355 15748 9411 15750
rect 10046 16088 10102 16144
rect 7483 15258 7539 15260
rect 7563 15258 7619 15260
rect 7643 15258 7699 15260
rect 7723 15258 7779 15260
rect 7483 15206 7529 15258
rect 7529 15206 7539 15258
rect 7563 15206 7593 15258
rect 7593 15206 7605 15258
rect 7605 15206 7619 15258
rect 7643 15206 7657 15258
rect 7657 15206 7669 15258
rect 7669 15206 7699 15258
rect 7723 15206 7733 15258
rect 7733 15206 7779 15258
rect 7483 15204 7539 15206
rect 7563 15204 7619 15206
rect 7643 15204 7699 15206
rect 7723 15204 7779 15206
rect 10046 15000 10102 15056
rect 9115 14714 9171 14716
rect 9195 14714 9251 14716
rect 9275 14714 9331 14716
rect 9355 14714 9411 14716
rect 9115 14662 9161 14714
rect 9161 14662 9171 14714
rect 9195 14662 9225 14714
rect 9225 14662 9237 14714
rect 9237 14662 9251 14714
rect 9275 14662 9289 14714
rect 9289 14662 9301 14714
rect 9301 14662 9331 14714
rect 9355 14662 9365 14714
rect 9365 14662 9411 14714
rect 9115 14660 9171 14662
rect 9195 14660 9251 14662
rect 9275 14660 9331 14662
rect 9355 14660 9411 14662
rect 7483 14170 7539 14172
rect 7563 14170 7619 14172
rect 7643 14170 7699 14172
rect 7723 14170 7779 14172
rect 7483 14118 7529 14170
rect 7529 14118 7539 14170
rect 7563 14118 7593 14170
rect 7593 14118 7605 14170
rect 7605 14118 7619 14170
rect 7643 14118 7657 14170
rect 7657 14118 7669 14170
rect 7669 14118 7699 14170
rect 7723 14118 7733 14170
rect 7733 14118 7779 14170
rect 7483 14116 7539 14118
rect 7563 14116 7619 14118
rect 7643 14116 7699 14118
rect 7723 14116 7779 14118
rect 10046 13912 10102 13968
rect 9115 13626 9171 13628
rect 9195 13626 9251 13628
rect 9275 13626 9331 13628
rect 9355 13626 9411 13628
rect 9115 13574 9161 13626
rect 9161 13574 9171 13626
rect 9195 13574 9225 13626
rect 9225 13574 9237 13626
rect 9237 13574 9251 13626
rect 9275 13574 9289 13626
rect 9289 13574 9301 13626
rect 9301 13574 9331 13626
rect 9355 13574 9365 13626
rect 9365 13574 9411 13626
rect 9115 13572 9171 13574
rect 9195 13572 9251 13574
rect 9275 13572 9331 13574
rect 9355 13572 9411 13574
rect 7483 13082 7539 13084
rect 7563 13082 7619 13084
rect 7643 13082 7699 13084
rect 7723 13082 7779 13084
rect 7483 13030 7529 13082
rect 7529 13030 7539 13082
rect 7563 13030 7593 13082
rect 7593 13030 7605 13082
rect 7605 13030 7619 13082
rect 7643 13030 7657 13082
rect 7657 13030 7669 13082
rect 7669 13030 7699 13082
rect 7723 13030 7733 13082
rect 7733 13030 7779 13082
rect 7483 13028 7539 13030
rect 7563 13028 7619 13030
rect 7643 13028 7699 13030
rect 7723 13028 7779 13030
rect 10046 12708 10102 12744
rect 10046 12688 10048 12708
rect 10048 12688 10100 12708
rect 10100 12688 10102 12708
rect 9115 12538 9171 12540
rect 9195 12538 9251 12540
rect 9275 12538 9331 12540
rect 9355 12538 9411 12540
rect 9115 12486 9161 12538
rect 9161 12486 9171 12538
rect 9195 12486 9225 12538
rect 9225 12486 9237 12538
rect 9237 12486 9251 12538
rect 9275 12486 9289 12538
rect 9289 12486 9301 12538
rect 9301 12486 9331 12538
rect 9355 12486 9365 12538
rect 9365 12486 9411 12538
rect 9115 12484 9171 12486
rect 9195 12484 9251 12486
rect 9275 12484 9331 12486
rect 9355 12484 9411 12486
rect 7483 11994 7539 11996
rect 7563 11994 7619 11996
rect 7643 11994 7699 11996
rect 7723 11994 7779 11996
rect 7483 11942 7529 11994
rect 7529 11942 7539 11994
rect 7563 11942 7593 11994
rect 7593 11942 7605 11994
rect 7605 11942 7619 11994
rect 7643 11942 7657 11994
rect 7657 11942 7669 11994
rect 7669 11942 7699 11994
rect 7723 11942 7733 11994
rect 7733 11942 7779 11994
rect 7483 11940 7539 11942
rect 7563 11940 7619 11942
rect 7643 11940 7699 11942
rect 7723 11940 7779 11942
rect 10046 11620 10102 11656
rect 10046 11600 10048 11620
rect 10048 11600 10100 11620
rect 10100 11600 10102 11620
rect 9115 11450 9171 11452
rect 9195 11450 9251 11452
rect 9275 11450 9331 11452
rect 9355 11450 9411 11452
rect 9115 11398 9161 11450
rect 9161 11398 9171 11450
rect 9195 11398 9225 11450
rect 9225 11398 9237 11450
rect 9237 11398 9251 11450
rect 9275 11398 9289 11450
rect 9289 11398 9301 11450
rect 9301 11398 9331 11450
rect 9355 11398 9365 11450
rect 9365 11398 9411 11450
rect 9115 11396 9171 11398
rect 9195 11396 9251 11398
rect 9275 11396 9331 11398
rect 9355 11396 9411 11398
rect 7483 10906 7539 10908
rect 7563 10906 7619 10908
rect 7643 10906 7699 10908
rect 7723 10906 7779 10908
rect 7483 10854 7529 10906
rect 7529 10854 7539 10906
rect 7563 10854 7593 10906
rect 7593 10854 7605 10906
rect 7605 10854 7619 10906
rect 7643 10854 7657 10906
rect 7657 10854 7669 10906
rect 7669 10854 7699 10906
rect 7723 10854 7733 10906
rect 7733 10854 7779 10906
rect 7483 10852 7539 10854
rect 7563 10852 7619 10854
rect 7643 10852 7699 10854
rect 7723 10852 7779 10854
rect 10046 10532 10102 10568
rect 10046 10512 10048 10532
rect 10048 10512 10100 10532
rect 10100 10512 10102 10532
rect 9115 10362 9171 10364
rect 9195 10362 9251 10364
rect 9275 10362 9331 10364
rect 9355 10362 9411 10364
rect 9115 10310 9161 10362
rect 9161 10310 9171 10362
rect 9195 10310 9225 10362
rect 9225 10310 9237 10362
rect 9237 10310 9251 10362
rect 9275 10310 9289 10362
rect 9289 10310 9301 10362
rect 9301 10310 9331 10362
rect 9355 10310 9365 10362
rect 9365 10310 9411 10362
rect 9115 10308 9171 10310
rect 9195 10308 9251 10310
rect 9275 10308 9331 10310
rect 9355 10308 9411 10310
rect 7483 9818 7539 9820
rect 7563 9818 7619 9820
rect 7643 9818 7699 9820
rect 7723 9818 7779 9820
rect 7483 9766 7529 9818
rect 7529 9766 7539 9818
rect 7563 9766 7593 9818
rect 7593 9766 7605 9818
rect 7605 9766 7619 9818
rect 7643 9766 7657 9818
rect 7657 9766 7669 9818
rect 7669 9766 7699 9818
rect 7723 9766 7733 9818
rect 7733 9766 7779 9818
rect 7483 9764 7539 9766
rect 7563 9764 7619 9766
rect 7643 9764 7699 9766
rect 7723 9764 7779 9766
rect 10046 9444 10102 9480
rect 10046 9424 10048 9444
rect 10048 9424 10100 9444
rect 10100 9424 10102 9444
rect 9115 9274 9171 9276
rect 9195 9274 9251 9276
rect 9275 9274 9331 9276
rect 9355 9274 9411 9276
rect 9115 9222 9161 9274
rect 9161 9222 9171 9274
rect 9195 9222 9225 9274
rect 9225 9222 9237 9274
rect 9237 9222 9251 9274
rect 9275 9222 9289 9274
rect 9289 9222 9301 9274
rect 9301 9222 9331 9274
rect 9355 9222 9365 9274
rect 9365 9222 9411 9274
rect 9115 9220 9171 9222
rect 9195 9220 9251 9222
rect 9275 9220 9331 9222
rect 9355 9220 9411 9222
rect 7483 8730 7539 8732
rect 7563 8730 7619 8732
rect 7643 8730 7699 8732
rect 7723 8730 7779 8732
rect 7483 8678 7529 8730
rect 7529 8678 7539 8730
rect 7563 8678 7593 8730
rect 7593 8678 7605 8730
rect 7605 8678 7619 8730
rect 7643 8678 7657 8730
rect 7657 8678 7669 8730
rect 7669 8678 7699 8730
rect 7723 8678 7733 8730
rect 7733 8678 7779 8730
rect 7483 8676 7539 8678
rect 7563 8676 7619 8678
rect 7643 8676 7699 8678
rect 7723 8676 7779 8678
rect 10046 8356 10102 8392
rect 10046 8336 10048 8356
rect 10048 8336 10100 8356
rect 10100 8336 10102 8356
rect 9115 8186 9171 8188
rect 9195 8186 9251 8188
rect 9275 8186 9331 8188
rect 9355 8186 9411 8188
rect 9115 8134 9161 8186
rect 9161 8134 9171 8186
rect 9195 8134 9225 8186
rect 9225 8134 9237 8186
rect 9237 8134 9251 8186
rect 9275 8134 9289 8186
rect 9289 8134 9301 8186
rect 9301 8134 9331 8186
rect 9355 8134 9365 8186
rect 9365 8134 9411 8186
rect 9115 8132 9171 8134
rect 9195 8132 9251 8134
rect 9275 8132 9331 8134
rect 9355 8132 9411 8134
rect 7483 7642 7539 7644
rect 7563 7642 7619 7644
rect 7643 7642 7699 7644
rect 7723 7642 7779 7644
rect 7483 7590 7529 7642
rect 7529 7590 7539 7642
rect 7563 7590 7593 7642
rect 7593 7590 7605 7642
rect 7605 7590 7619 7642
rect 7643 7590 7657 7642
rect 7657 7590 7669 7642
rect 7669 7590 7699 7642
rect 7723 7590 7733 7642
rect 7733 7590 7779 7642
rect 7483 7588 7539 7590
rect 7563 7588 7619 7590
rect 7643 7588 7699 7590
rect 7723 7588 7779 7590
rect 10046 7268 10102 7304
rect 10046 7248 10048 7268
rect 10048 7248 10100 7268
rect 10100 7248 10102 7268
rect 9115 7098 9171 7100
rect 9195 7098 9251 7100
rect 9275 7098 9331 7100
rect 9355 7098 9411 7100
rect 9115 7046 9161 7098
rect 9161 7046 9171 7098
rect 9195 7046 9225 7098
rect 9225 7046 9237 7098
rect 9237 7046 9251 7098
rect 9275 7046 9289 7098
rect 9289 7046 9301 7098
rect 9301 7046 9331 7098
rect 9355 7046 9365 7098
rect 9365 7046 9411 7098
rect 9115 7044 9171 7046
rect 9195 7044 9251 7046
rect 9275 7044 9331 7046
rect 9355 7044 9411 7046
rect 7483 6554 7539 6556
rect 7563 6554 7619 6556
rect 7643 6554 7699 6556
rect 7723 6554 7779 6556
rect 7483 6502 7529 6554
rect 7529 6502 7539 6554
rect 7563 6502 7593 6554
rect 7593 6502 7605 6554
rect 7605 6502 7619 6554
rect 7643 6502 7657 6554
rect 7657 6502 7669 6554
rect 7669 6502 7699 6554
rect 7723 6502 7733 6554
rect 7733 6502 7779 6554
rect 7483 6500 7539 6502
rect 7563 6500 7619 6502
rect 7643 6500 7699 6502
rect 7723 6500 7779 6502
rect 10046 6060 10048 6080
rect 10048 6060 10100 6080
rect 10100 6060 10102 6080
rect 5851 6010 5907 6012
rect 5931 6010 5987 6012
rect 6011 6010 6067 6012
rect 6091 6010 6147 6012
rect 5851 5958 5897 6010
rect 5897 5958 5907 6010
rect 5931 5958 5961 6010
rect 5961 5958 5973 6010
rect 5973 5958 5987 6010
rect 6011 5958 6025 6010
rect 6025 5958 6037 6010
rect 6037 5958 6067 6010
rect 6091 5958 6101 6010
rect 6101 5958 6147 6010
rect 5851 5956 5907 5958
rect 5931 5956 5987 5958
rect 6011 5956 6067 5958
rect 6091 5956 6147 5958
rect 9115 6010 9171 6012
rect 9195 6010 9251 6012
rect 9275 6010 9331 6012
rect 9355 6010 9411 6012
rect 9115 5958 9161 6010
rect 9161 5958 9171 6010
rect 9195 5958 9225 6010
rect 9225 5958 9237 6010
rect 9237 5958 9251 6010
rect 9275 5958 9289 6010
rect 9289 5958 9301 6010
rect 9301 5958 9331 6010
rect 9355 5958 9365 6010
rect 9365 5958 9411 6010
rect 9115 5956 9171 5958
rect 9195 5956 9251 5958
rect 9275 5956 9331 5958
rect 9355 5956 9411 5958
rect 4219 5466 4275 5468
rect 4299 5466 4355 5468
rect 4379 5466 4435 5468
rect 4459 5466 4515 5468
rect 4219 5414 4265 5466
rect 4265 5414 4275 5466
rect 4299 5414 4329 5466
rect 4329 5414 4341 5466
rect 4341 5414 4355 5466
rect 4379 5414 4393 5466
rect 4393 5414 4405 5466
rect 4405 5414 4435 5466
rect 4459 5414 4469 5466
rect 4469 5414 4515 5466
rect 4219 5412 4275 5414
rect 4299 5412 4355 5414
rect 4379 5412 4435 5414
rect 4459 5412 4515 5414
rect 7483 5466 7539 5468
rect 7563 5466 7619 5468
rect 7643 5466 7699 5468
rect 7723 5466 7779 5468
rect 7483 5414 7529 5466
rect 7529 5414 7539 5466
rect 7563 5414 7593 5466
rect 7593 5414 7605 5466
rect 7605 5414 7619 5466
rect 7643 5414 7657 5466
rect 7657 5414 7669 5466
rect 7669 5414 7699 5466
rect 7723 5414 7733 5466
rect 7733 5414 7779 5466
rect 7483 5412 7539 5414
rect 7563 5412 7619 5414
rect 7643 5412 7699 5414
rect 7723 5412 7779 5414
rect 10046 6024 10102 6060
rect 4219 4378 4275 4380
rect 4299 4378 4355 4380
rect 4379 4378 4435 4380
rect 4459 4378 4515 4380
rect 4219 4326 4265 4378
rect 4265 4326 4275 4378
rect 4299 4326 4329 4378
rect 4329 4326 4341 4378
rect 4341 4326 4355 4378
rect 4379 4326 4393 4378
rect 4393 4326 4405 4378
rect 4405 4326 4435 4378
rect 4459 4326 4469 4378
rect 4469 4326 4515 4378
rect 4219 4324 4275 4326
rect 4299 4324 4355 4326
rect 4379 4324 4435 4326
rect 4459 4324 4515 4326
rect 5851 4922 5907 4924
rect 5931 4922 5987 4924
rect 6011 4922 6067 4924
rect 6091 4922 6147 4924
rect 5851 4870 5897 4922
rect 5897 4870 5907 4922
rect 5931 4870 5961 4922
rect 5961 4870 5973 4922
rect 5973 4870 5987 4922
rect 6011 4870 6025 4922
rect 6025 4870 6037 4922
rect 6037 4870 6067 4922
rect 6091 4870 6101 4922
rect 6101 4870 6147 4922
rect 5851 4868 5907 4870
rect 5931 4868 5987 4870
rect 6011 4868 6067 4870
rect 6091 4868 6147 4870
rect 9115 4922 9171 4924
rect 9195 4922 9251 4924
rect 9275 4922 9331 4924
rect 9355 4922 9411 4924
rect 9115 4870 9161 4922
rect 9161 4870 9171 4922
rect 9195 4870 9225 4922
rect 9225 4870 9237 4922
rect 9237 4870 9251 4922
rect 9275 4870 9289 4922
rect 9289 4870 9301 4922
rect 9301 4870 9331 4922
rect 9355 4870 9365 4922
rect 9365 4870 9411 4922
rect 9115 4868 9171 4870
rect 9195 4868 9251 4870
rect 9275 4868 9331 4870
rect 9355 4868 9411 4870
rect 7483 4378 7539 4380
rect 7563 4378 7619 4380
rect 7643 4378 7699 4380
rect 7723 4378 7779 4380
rect 7483 4326 7529 4378
rect 7529 4326 7539 4378
rect 7563 4326 7593 4378
rect 7593 4326 7605 4378
rect 7605 4326 7619 4378
rect 7643 4326 7657 4378
rect 7657 4326 7669 4378
rect 7669 4326 7699 4378
rect 7723 4326 7733 4378
rect 7733 4326 7779 4378
rect 7483 4324 7539 4326
rect 7563 4324 7619 4326
rect 7643 4324 7699 4326
rect 7723 4324 7779 4326
rect 5851 3834 5907 3836
rect 5931 3834 5987 3836
rect 6011 3834 6067 3836
rect 6091 3834 6147 3836
rect 5851 3782 5897 3834
rect 5897 3782 5907 3834
rect 5931 3782 5961 3834
rect 5961 3782 5973 3834
rect 5973 3782 5987 3834
rect 6011 3782 6025 3834
rect 6025 3782 6037 3834
rect 6037 3782 6067 3834
rect 6091 3782 6101 3834
rect 6101 3782 6147 3834
rect 5851 3780 5907 3782
rect 5931 3780 5987 3782
rect 6011 3780 6067 3782
rect 6091 3780 6147 3782
rect 9115 3834 9171 3836
rect 9195 3834 9251 3836
rect 9275 3834 9331 3836
rect 9355 3834 9411 3836
rect 9115 3782 9161 3834
rect 9161 3782 9171 3834
rect 9195 3782 9225 3834
rect 9225 3782 9237 3834
rect 9237 3782 9251 3834
rect 9275 3782 9289 3834
rect 9289 3782 9301 3834
rect 9301 3782 9331 3834
rect 9355 3782 9365 3834
rect 9365 3782 9411 3834
rect 9115 3780 9171 3782
rect 9195 3780 9251 3782
rect 9275 3780 9331 3782
rect 9355 3780 9411 3782
rect 10046 4972 10048 4992
rect 10048 4972 10100 4992
rect 10100 4972 10102 4992
rect 10046 4936 10102 4972
rect 10046 3884 10048 3904
rect 10048 3884 10100 3904
rect 10100 3884 10102 3904
rect 10046 3848 10102 3884
rect 4219 3290 4275 3292
rect 4299 3290 4355 3292
rect 4379 3290 4435 3292
rect 4459 3290 4515 3292
rect 4219 3238 4265 3290
rect 4265 3238 4275 3290
rect 4299 3238 4329 3290
rect 4329 3238 4341 3290
rect 4341 3238 4355 3290
rect 4379 3238 4393 3290
rect 4393 3238 4405 3290
rect 4405 3238 4435 3290
rect 4459 3238 4469 3290
rect 4469 3238 4515 3290
rect 4219 3236 4275 3238
rect 4299 3236 4355 3238
rect 4379 3236 4435 3238
rect 4459 3236 4515 3238
rect 7483 3290 7539 3292
rect 7563 3290 7619 3292
rect 7643 3290 7699 3292
rect 7723 3290 7779 3292
rect 7483 3238 7529 3290
rect 7529 3238 7539 3290
rect 7563 3238 7593 3290
rect 7593 3238 7605 3290
rect 7605 3238 7619 3290
rect 7643 3238 7657 3290
rect 7657 3238 7669 3290
rect 7669 3238 7699 3290
rect 7723 3238 7733 3290
rect 7733 3238 7779 3290
rect 7483 3236 7539 3238
rect 7563 3236 7619 3238
rect 7643 3236 7699 3238
rect 7723 3236 7779 3238
rect 2588 2746 2644 2748
rect 2668 2746 2724 2748
rect 2748 2746 2804 2748
rect 2828 2746 2884 2748
rect 2588 2694 2634 2746
rect 2634 2694 2644 2746
rect 2668 2694 2698 2746
rect 2698 2694 2710 2746
rect 2710 2694 2724 2746
rect 2748 2694 2762 2746
rect 2762 2694 2774 2746
rect 2774 2694 2804 2746
rect 2828 2694 2838 2746
rect 2838 2694 2884 2746
rect 2588 2692 2644 2694
rect 2668 2692 2724 2694
rect 2748 2692 2804 2694
rect 2828 2692 2884 2694
rect 5851 2746 5907 2748
rect 5931 2746 5987 2748
rect 6011 2746 6067 2748
rect 6091 2746 6147 2748
rect 5851 2694 5897 2746
rect 5897 2694 5907 2746
rect 5931 2694 5961 2746
rect 5961 2694 5973 2746
rect 5973 2694 5987 2746
rect 6011 2694 6025 2746
rect 6025 2694 6037 2746
rect 6037 2694 6067 2746
rect 6091 2694 6101 2746
rect 6101 2694 6147 2746
rect 5851 2692 5907 2694
rect 5931 2692 5987 2694
rect 6011 2692 6067 2694
rect 6091 2692 6147 2694
rect 10046 2760 10102 2816
rect 9115 2746 9171 2748
rect 9195 2746 9251 2748
rect 9275 2746 9331 2748
rect 9355 2746 9411 2748
rect 9115 2694 9161 2746
rect 9161 2694 9171 2746
rect 9195 2694 9225 2746
rect 9225 2694 9237 2746
rect 9237 2694 9251 2746
rect 9275 2694 9289 2746
rect 9289 2694 9301 2746
rect 9301 2694 9331 2746
rect 9355 2694 9365 2746
rect 9365 2694 9411 2746
rect 9115 2692 9171 2694
rect 9195 2692 9251 2694
rect 9275 2692 9331 2694
rect 9355 2692 9411 2694
rect 1398 2352 1454 2408
rect 1306 1400 1362 1456
rect 4219 2202 4275 2204
rect 4299 2202 4355 2204
rect 4379 2202 4435 2204
rect 4459 2202 4515 2204
rect 4219 2150 4265 2202
rect 4265 2150 4275 2202
rect 4299 2150 4329 2202
rect 4329 2150 4341 2202
rect 4341 2150 4355 2202
rect 4379 2150 4393 2202
rect 4393 2150 4405 2202
rect 4405 2150 4435 2202
rect 4459 2150 4469 2202
rect 4469 2150 4515 2202
rect 4219 2148 4275 2150
rect 4299 2148 4355 2150
rect 4379 2148 4435 2150
rect 4459 2148 4515 2150
rect 7483 2202 7539 2204
rect 7563 2202 7619 2204
rect 7643 2202 7699 2204
rect 7723 2202 7779 2204
rect 7483 2150 7529 2202
rect 7529 2150 7539 2202
rect 7563 2150 7593 2202
rect 7593 2150 7605 2202
rect 7605 2150 7619 2202
rect 7643 2150 7657 2202
rect 7657 2150 7669 2202
rect 7669 2150 7699 2202
rect 7723 2150 7733 2202
rect 7733 2150 7779 2202
rect 7483 2148 7539 2150
rect 7563 2148 7619 2150
rect 7643 2148 7699 2150
rect 7723 2148 7779 2150
rect 2778 1944 2834 2000
rect 10046 1672 10102 1728
rect 2042 992 2098 1048
rect 10966 620 10968 640
rect 10968 620 11020 640
rect 11020 620 11022 640
rect 10966 584 11022 620
<< metal3 >>
rect 0 79658 800 79688
rect 3141 79658 3207 79661
rect 0 79656 3207 79658
rect 0 79600 3146 79656
rect 3202 79600 3207 79656
rect 0 79598 3207 79600
rect 0 79568 800 79598
rect 3141 79595 3207 79598
rect 9489 79386 9555 79389
rect 11200 79386 12000 79416
rect 9489 79384 12000 79386
rect 9489 79328 9494 79384
rect 9550 79328 12000 79384
rect 9489 79326 12000 79328
rect 9489 79323 9555 79326
rect 11200 79296 12000 79326
rect 0 79250 800 79280
rect 3049 79250 3115 79253
rect 0 79248 3115 79250
rect 0 79192 3054 79248
rect 3110 79192 3115 79248
rect 0 79190 3115 79192
rect 0 79160 800 79190
rect 3049 79187 3115 79190
rect 0 78842 800 78872
rect 3969 78842 4035 78845
rect 0 78840 4035 78842
rect 0 78784 3974 78840
rect 4030 78784 4035 78840
rect 0 78782 4035 78784
rect 0 78752 800 78782
rect 3969 78779 4035 78782
rect 0 78298 800 78328
rect 2957 78298 3023 78301
rect 0 78296 3023 78298
rect 0 78240 2962 78296
rect 3018 78240 3023 78296
rect 0 78238 3023 78240
rect 0 78208 800 78238
rect 2957 78235 3023 78238
rect 10961 78298 11027 78301
rect 11200 78298 12000 78328
rect 10961 78296 12000 78298
rect 10961 78240 10966 78296
rect 11022 78240 12000 78296
rect 10961 78238 12000 78240
rect 10961 78235 11027 78238
rect 11200 78208 12000 78238
rect 0 77890 800 77920
rect 0 77830 1410 77890
rect 0 77800 800 77830
rect 1350 77618 1410 77830
rect 2576 77824 2896 77825
rect 2576 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2576 77759 2896 77760
rect 5839 77824 6159 77825
rect 5839 77760 5847 77824
rect 5911 77760 5927 77824
rect 5991 77760 6007 77824
rect 6071 77760 6087 77824
rect 6151 77760 6159 77824
rect 5839 77759 6159 77760
rect 9103 77824 9423 77825
rect 9103 77760 9111 77824
rect 9175 77760 9191 77824
rect 9255 77760 9271 77824
rect 9335 77760 9351 77824
rect 9415 77760 9423 77824
rect 9103 77759 9423 77760
rect 2865 77618 2931 77621
rect 1350 77616 2931 77618
rect 1350 77560 2870 77616
rect 2926 77560 2931 77616
rect 1350 77558 2931 77560
rect 2865 77555 2931 77558
rect 0 77482 800 77512
rect 2037 77482 2103 77485
rect 0 77480 2103 77482
rect 0 77424 2042 77480
rect 2098 77424 2103 77480
rect 0 77422 2103 77424
rect 0 77392 800 77422
rect 2037 77419 2103 77422
rect 4207 77280 4527 77281
rect 4207 77216 4215 77280
rect 4279 77216 4295 77280
rect 4359 77216 4375 77280
rect 4439 77216 4455 77280
rect 4519 77216 4527 77280
rect 4207 77215 4527 77216
rect 7471 77280 7791 77281
rect 7471 77216 7479 77280
rect 7543 77216 7559 77280
rect 7623 77216 7639 77280
rect 7703 77216 7719 77280
rect 7783 77216 7791 77280
rect 7471 77215 7791 77216
rect 10133 77210 10199 77213
rect 11200 77210 12000 77240
rect 10133 77208 12000 77210
rect 10133 77152 10138 77208
rect 10194 77152 12000 77208
rect 10133 77150 12000 77152
rect 10133 77147 10199 77150
rect 11200 77120 12000 77150
rect 0 76938 800 76968
rect 2037 76938 2103 76941
rect 0 76936 2103 76938
rect 0 76880 2042 76936
rect 2098 76880 2103 76936
rect 0 76878 2103 76880
rect 0 76848 800 76878
rect 2037 76875 2103 76878
rect 2576 76736 2896 76737
rect 2576 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2576 76671 2896 76672
rect 5839 76736 6159 76737
rect 5839 76672 5847 76736
rect 5911 76672 5927 76736
rect 5991 76672 6007 76736
rect 6071 76672 6087 76736
rect 6151 76672 6159 76736
rect 5839 76671 6159 76672
rect 9103 76736 9423 76737
rect 9103 76672 9111 76736
rect 9175 76672 9191 76736
rect 9255 76672 9271 76736
rect 9335 76672 9351 76736
rect 9415 76672 9423 76736
rect 9103 76671 9423 76672
rect 0 76530 800 76560
rect 1485 76530 1551 76533
rect 0 76528 1551 76530
rect 0 76472 1490 76528
rect 1546 76472 1551 76528
rect 0 76470 1551 76472
rect 0 76440 800 76470
rect 1485 76467 1551 76470
rect 4207 76192 4527 76193
rect 0 76122 800 76152
rect 4207 76128 4215 76192
rect 4279 76128 4295 76192
rect 4359 76128 4375 76192
rect 4439 76128 4455 76192
rect 4519 76128 4527 76192
rect 4207 76127 4527 76128
rect 7471 76192 7791 76193
rect 7471 76128 7479 76192
rect 7543 76128 7559 76192
rect 7623 76128 7639 76192
rect 7703 76128 7719 76192
rect 7783 76128 7791 76192
rect 7471 76127 7791 76128
rect 1393 76122 1459 76125
rect 0 76120 1459 76122
rect 0 76064 1398 76120
rect 1454 76064 1459 76120
rect 0 76062 1459 76064
rect 0 76032 800 76062
rect 1393 76059 1459 76062
rect 10133 76122 10199 76125
rect 11200 76122 12000 76152
rect 10133 76120 12000 76122
rect 10133 76064 10138 76120
rect 10194 76064 12000 76120
rect 10133 76062 12000 76064
rect 10133 76059 10199 76062
rect 11200 76032 12000 76062
rect 2576 75648 2896 75649
rect 0 75578 800 75608
rect 2576 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2576 75583 2896 75584
rect 5839 75648 6159 75649
rect 5839 75584 5847 75648
rect 5911 75584 5927 75648
rect 5991 75584 6007 75648
rect 6071 75584 6087 75648
rect 6151 75584 6159 75648
rect 5839 75583 6159 75584
rect 9103 75648 9423 75649
rect 9103 75584 9111 75648
rect 9175 75584 9191 75648
rect 9255 75584 9271 75648
rect 9335 75584 9351 75648
rect 9415 75584 9423 75648
rect 9103 75583 9423 75584
rect 2221 75578 2287 75581
rect 0 75576 2287 75578
rect 0 75520 2226 75576
rect 2282 75520 2287 75576
rect 0 75518 2287 75520
rect 0 75488 800 75518
rect 2221 75515 2287 75518
rect 0 75170 800 75200
rect 1301 75170 1367 75173
rect 0 75168 1367 75170
rect 0 75112 1306 75168
rect 1362 75112 1367 75168
rect 0 75110 1367 75112
rect 0 75080 800 75110
rect 1301 75107 1367 75110
rect 4207 75104 4527 75105
rect 4207 75040 4215 75104
rect 4279 75040 4295 75104
rect 4359 75040 4375 75104
rect 4439 75040 4455 75104
rect 4519 75040 4527 75104
rect 4207 75039 4527 75040
rect 7471 75104 7791 75105
rect 7471 75040 7479 75104
rect 7543 75040 7559 75104
rect 7623 75040 7639 75104
rect 7703 75040 7719 75104
rect 7783 75040 7791 75104
rect 7471 75039 7791 75040
rect 10133 75034 10199 75037
rect 11200 75034 12000 75064
rect 10133 75032 12000 75034
rect 10133 74976 10138 75032
rect 10194 74976 12000 75032
rect 10133 74974 12000 74976
rect 10133 74971 10199 74974
rect 11200 74944 12000 74974
rect 0 74762 800 74792
rect 2773 74762 2839 74765
rect 0 74760 2839 74762
rect 0 74704 2778 74760
rect 2834 74704 2839 74760
rect 0 74702 2839 74704
rect 0 74672 800 74702
rect 2773 74699 2839 74702
rect 2576 74560 2896 74561
rect 2576 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2576 74495 2896 74496
rect 5839 74560 6159 74561
rect 5839 74496 5847 74560
rect 5911 74496 5927 74560
rect 5991 74496 6007 74560
rect 6071 74496 6087 74560
rect 6151 74496 6159 74560
rect 5839 74495 6159 74496
rect 9103 74560 9423 74561
rect 9103 74496 9111 74560
rect 9175 74496 9191 74560
rect 9255 74496 9271 74560
rect 9335 74496 9351 74560
rect 9415 74496 9423 74560
rect 9103 74495 9423 74496
rect 0 74354 800 74384
rect 1393 74354 1459 74357
rect 0 74352 1459 74354
rect 0 74296 1398 74352
rect 1454 74296 1459 74352
rect 0 74294 1459 74296
rect 0 74264 800 74294
rect 1393 74291 1459 74294
rect 4207 74016 4527 74017
rect 4207 73952 4215 74016
rect 4279 73952 4295 74016
rect 4359 73952 4375 74016
rect 4439 73952 4455 74016
rect 4519 73952 4527 74016
rect 4207 73951 4527 73952
rect 7471 74016 7791 74017
rect 7471 73952 7479 74016
rect 7543 73952 7559 74016
rect 7623 73952 7639 74016
rect 7703 73952 7719 74016
rect 7783 73952 7791 74016
rect 7471 73951 7791 73952
rect 10133 73946 10199 73949
rect 11200 73946 12000 73976
rect 10133 73944 12000 73946
rect 10133 73888 10138 73944
rect 10194 73888 12000 73944
rect 10133 73886 12000 73888
rect 10133 73883 10199 73886
rect 11200 73856 12000 73886
rect 0 73810 800 73840
rect 2865 73810 2931 73813
rect 0 73808 2931 73810
rect 0 73752 2870 73808
rect 2926 73752 2931 73808
rect 0 73750 2931 73752
rect 0 73720 800 73750
rect 2865 73747 2931 73750
rect 2576 73472 2896 73473
rect 0 73402 800 73432
rect 2576 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2576 73407 2896 73408
rect 5839 73472 6159 73473
rect 5839 73408 5847 73472
rect 5911 73408 5927 73472
rect 5991 73408 6007 73472
rect 6071 73408 6087 73472
rect 6151 73408 6159 73472
rect 5839 73407 6159 73408
rect 9103 73472 9423 73473
rect 9103 73408 9111 73472
rect 9175 73408 9191 73472
rect 9255 73408 9271 73472
rect 9335 73408 9351 73472
rect 9415 73408 9423 73472
rect 9103 73407 9423 73408
rect 1301 73402 1367 73405
rect 0 73400 1367 73402
rect 0 73344 1306 73400
rect 1362 73344 1367 73400
rect 0 73342 1367 73344
rect 0 73312 800 73342
rect 1301 73339 1367 73342
rect 0 72994 800 73024
rect 1393 72994 1459 72997
rect 0 72992 1459 72994
rect 0 72936 1398 72992
rect 1454 72936 1459 72992
rect 0 72934 1459 72936
rect 0 72904 800 72934
rect 1393 72931 1459 72934
rect 4207 72928 4527 72929
rect 4207 72864 4215 72928
rect 4279 72864 4295 72928
rect 4359 72864 4375 72928
rect 4439 72864 4455 72928
rect 4519 72864 4527 72928
rect 4207 72863 4527 72864
rect 7471 72928 7791 72929
rect 7471 72864 7479 72928
rect 7543 72864 7559 72928
rect 7623 72864 7639 72928
rect 7703 72864 7719 72928
rect 7783 72864 7791 72928
rect 7471 72863 7791 72864
rect 10133 72722 10199 72725
rect 11200 72722 12000 72752
rect 10133 72720 12000 72722
rect 10133 72664 10138 72720
rect 10194 72664 12000 72720
rect 10133 72662 12000 72664
rect 10133 72659 10199 72662
rect 11200 72632 12000 72662
rect 0 72450 800 72480
rect 2037 72450 2103 72453
rect 0 72448 2103 72450
rect 0 72392 2042 72448
rect 2098 72392 2103 72448
rect 0 72390 2103 72392
rect 0 72360 800 72390
rect 2037 72387 2103 72390
rect 2576 72384 2896 72385
rect 2576 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2576 72319 2896 72320
rect 5839 72384 6159 72385
rect 5839 72320 5847 72384
rect 5911 72320 5927 72384
rect 5991 72320 6007 72384
rect 6071 72320 6087 72384
rect 6151 72320 6159 72384
rect 5839 72319 6159 72320
rect 9103 72384 9423 72385
rect 9103 72320 9111 72384
rect 9175 72320 9191 72384
rect 9255 72320 9271 72384
rect 9335 72320 9351 72384
rect 9415 72320 9423 72384
rect 9103 72319 9423 72320
rect 0 72042 800 72072
rect 1301 72042 1367 72045
rect 0 72040 1367 72042
rect 0 71984 1306 72040
rect 1362 71984 1367 72040
rect 0 71982 1367 71984
rect 0 71952 800 71982
rect 1301 71979 1367 71982
rect 4207 71840 4527 71841
rect 4207 71776 4215 71840
rect 4279 71776 4295 71840
rect 4359 71776 4375 71840
rect 4439 71776 4455 71840
rect 4519 71776 4527 71840
rect 4207 71775 4527 71776
rect 7471 71840 7791 71841
rect 7471 71776 7479 71840
rect 7543 71776 7559 71840
rect 7623 71776 7639 71840
rect 7703 71776 7719 71840
rect 7783 71776 7791 71840
rect 7471 71775 7791 71776
rect 0 71634 800 71664
rect 1209 71634 1275 71637
rect 0 71632 1275 71634
rect 0 71576 1214 71632
rect 1270 71576 1275 71632
rect 0 71574 1275 71576
rect 0 71544 800 71574
rect 1209 71571 1275 71574
rect 10133 71634 10199 71637
rect 11200 71634 12000 71664
rect 10133 71632 12000 71634
rect 10133 71576 10138 71632
rect 10194 71576 12000 71632
rect 10133 71574 12000 71576
rect 10133 71571 10199 71574
rect 11200 71544 12000 71574
rect 2576 71296 2896 71297
rect 2576 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2576 71231 2896 71232
rect 5839 71296 6159 71297
rect 5839 71232 5847 71296
rect 5911 71232 5927 71296
rect 5991 71232 6007 71296
rect 6071 71232 6087 71296
rect 6151 71232 6159 71296
rect 5839 71231 6159 71232
rect 9103 71296 9423 71297
rect 9103 71232 9111 71296
rect 9175 71232 9191 71296
rect 9255 71232 9271 71296
rect 9335 71232 9351 71296
rect 9415 71232 9423 71296
rect 9103 71231 9423 71232
rect 0 71090 800 71120
rect 1393 71090 1459 71093
rect 0 71088 1459 71090
rect 0 71032 1398 71088
rect 1454 71032 1459 71088
rect 0 71030 1459 71032
rect 0 71000 800 71030
rect 1393 71027 1459 71030
rect 4207 70752 4527 70753
rect 0 70682 800 70712
rect 4207 70688 4215 70752
rect 4279 70688 4295 70752
rect 4359 70688 4375 70752
rect 4439 70688 4455 70752
rect 4519 70688 4527 70752
rect 4207 70687 4527 70688
rect 7471 70752 7791 70753
rect 7471 70688 7479 70752
rect 7543 70688 7559 70752
rect 7623 70688 7639 70752
rect 7703 70688 7719 70752
rect 7783 70688 7791 70752
rect 7471 70687 7791 70688
rect 2773 70682 2839 70685
rect 0 70680 2839 70682
rect 0 70624 2778 70680
rect 2834 70624 2839 70680
rect 0 70622 2839 70624
rect 0 70592 800 70622
rect 2773 70619 2839 70622
rect 1526 70484 1532 70548
rect 1596 70546 1602 70548
rect 1669 70546 1735 70549
rect 1596 70544 1735 70546
rect 1596 70488 1674 70544
rect 1730 70488 1735 70544
rect 1596 70486 1735 70488
rect 1596 70484 1602 70486
rect 1669 70483 1735 70486
rect 10133 70546 10199 70549
rect 11200 70546 12000 70576
rect 10133 70544 12000 70546
rect 10133 70488 10138 70544
rect 10194 70488 12000 70544
rect 10133 70486 12000 70488
rect 10133 70483 10199 70486
rect 11200 70456 12000 70486
rect 0 70274 800 70304
rect 1301 70274 1367 70277
rect 0 70272 1367 70274
rect 0 70216 1306 70272
rect 1362 70216 1367 70272
rect 0 70214 1367 70216
rect 0 70184 800 70214
rect 1301 70211 1367 70214
rect 2576 70208 2896 70209
rect 2576 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2576 70143 2896 70144
rect 5839 70208 6159 70209
rect 5839 70144 5847 70208
rect 5911 70144 5927 70208
rect 5991 70144 6007 70208
rect 6071 70144 6087 70208
rect 6151 70144 6159 70208
rect 5839 70143 6159 70144
rect 9103 70208 9423 70209
rect 9103 70144 9111 70208
rect 9175 70144 9191 70208
rect 9255 70144 9271 70208
rect 9335 70144 9351 70208
rect 9415 70144 9423 70208
rect 9103 70143 9423 70144
rect 0 69866 800 69896
rect 2865 69866 2931 69869
rect 0 69864 2931 69866
rect 0 69808 2870 69864
rect 2926 69808 2931 69864
rect 0 69806 2931 69808
rect 0 69776 800 69806
rect 2865 69803 2931 69806
rect 4207 69664 4527 69665
rect 4207 69600 4215 69664
rect 4279 69600 4295 69664
rect 4359 69600 4375 69664
rect 4439 69600 4455 69664
rect 4519 69600 4527 69664
rect 4207 69599 4527 69600
rect 7471 69664 7791 69665
rect 7471 69600 7479 69664
rect 7543 69600 7559 69664
rect 7623 69600 7639 69664
rect 7703 69600 7719 69664
rect 7783 69600 7791 69664
rect 7471 69599 7791 69600
rect 10133 69458 10199 69461
rect 11200 69458 12000 69488
rect 10133 69456 12000 69458
rect 10133 69400 10138 69456
rect 10194 69400 12000 69456
rect 10133 69398 12000 69400
rect 10133 69395 10199 69398
rect 11200 69368 12000 69398
rect 0 69322 800 69352
rect 1209 69322 1275 69325
rect 0 69320 1275 69322
rect 0 69264 1214 69320
rect 1270 69264 1275 69320
rect 0 69262 1275 69264
rect 0 69232 800 69262
rect 1209 69259 1275 69262
rect 2576 69120 2896 69121
rect 2576 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2576 69055 2896 69056
rect 5839 69120 6159 69121
rect 5839 69056 5847 69120
rect 5911 69056 5927 69120
rect 5991 69056 6007 69120
rect 6071 69056 6087 69120
rect 6151 69056 6159 69120
rect 5839 69055 6159 69056
rect 9103 69120 9423 69121
rect 9103 69056 9111 69120
rect 9175 69056 9191 69120
rect 9255 69056 9271 69120
rect 9335 69056 9351 69120
rect 9415 69056 9423 69120
rect 9103 69055 9423 69056
rect 1710 68988 1716 69052
rect 1780 69050 1786 69052
rect 2313 69050 2379 69053
rect 1780 69048 2379 69050
rect 1780 68992 2318 69048
rect 2374 68992 2379 69048
rect 1780 68990 2379 68992
rect 1780 68988 1786 68990
rect 2313 68987 2379 68990
rect 0 68914 800 68944
rect 1393 68914 1459 68917
rect 0 68912 1459 68914
rect 0 68856 1398 68912
rect 1454 68856 1459 68912
rect 0 68854 1459 68856
rect 0 68824 800 68854
rect 1393 68851 1459 68854
rect 2078 68580 2084 68644
rect 2148 68642 2154 68644
rect 2221 68642 2287 68645
rect 2148 68640 2287 68642
rect 2148 68584 2226 68640
rect 2282 68584 2287 68640
rect 2148 68582 2287 68584
rect 2148 68580 2154 68582
rect 2221 68579 2287 68582
rect 4207 68576 4527 68577
rect 0 68506 800 68536
rect 4207 68512 4215 68576
rect 4279 68512 4295 68576
rect 4359 68512 4375 68576
rect 4439 68512 4455 68576
rect 4519 68512 4527 68576
rect 4207 68511 4527 68512
rect 7471 68576 7791 68577
rect 7471 68512 7479 68576
rect 7543 68512 7559 68576
rect 7623 68512 7639 68576
rect 7703 68512 7719 68576
rect 7783 68512 7791 68576
rect 7471 68511 7791 68512
rect 1301 68506 1367 68509
rect 0 68504 1367 68506
rect 0 68448 1306 68504
rect 1362 68448 1367 68504
rect 0 68446 1367 68448
rect 0 68416 800 68446
rect 1301 68443 1367 68446
rect 10133 68370 10199 68373
rect 11200 68370 12000 68400
rect 10133 68368 12000 68370
rect 10133 68312 10138 68368
rect 10194 68312 12000 68368
rect 10133 68310 12000 68312
rect 10133 68307 10199 68310
rect 11200 68280 12000 68310
rect 2576 68032 2896 68033
rect 0 67962 800 67992
rect 2576 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2576 67967 2896 67968
rect 5839 68032 6159 68033
rect 5839 67968 5847 68032
rect 5911 67968 5927 68032
rect 5991 67968 6007 68032
rect 6071 67968 6087 68032
rect 6151 67968 6159 68032
rect 5839 67967 6159 67968
rect 9103 68032 9423 68033
rect 9103 67968 9111 68032
rect 9175 67968 9191 68032
rect 9255 67968 9271 68032
rect 9335 67968 9351 68032
rect 9415 67968 9423 68032
rect 9103 67967 9423 67968
rect 1393 67962 1459 67965
rect 0 67960 1459 67962
rect 0 67904 1398 67960
rect 1454 67904 1459 67960
rect 0 67902 1459 67904
rect 0 67872 800 67902
rect 1393 67899 1459 67902
rect 1485 67828 1551 67829
rect 1485 67824 1532 67828
rect 1596 67826 1602 67828
rect 1485 67768 1490 67824
rect 1485 67764 1532 67768
rect 1596 67766 1642 67826
rect 1596 67764 1602 67766
rect 1485 67763 1551 67764
rect 0 67554 800 67584
rect 1393 67554 1459 67557
rect 0 67552 1459 67554
rect 0 67496 1398 67552
rect 1454 67496 1459 67552
rect 0 67494 1459 67496
rect 0 67464 800 67494
rect 1393 67491 1459 67494
rect 4207 67488 4527 67489
rect 4207 67424 4215 67488
rect 4279 67424 4295 67488
rect 4359 67424 4375 67488
rect 4439 67424 4455 67488
rect 4519 67424 4527 67488
rect 4207 67423 4527 67424
rect 7471 67488 7791 67489
rect 7471 67424 7479 67488
rect 7543 67424 7559 67488
rect 7623 67424 7639 67488
rect 7703 67424 7719 67488
rect 7783 67424 7791 67488
rect 7471 67423 7791 67424
rect 10133 67282 10199 67285
rect 11200 67282 12000 67312
rect 10133 67280 12000 67282
rect 10133 67224 10138 67280
rect 10194 67224 12000 67280
rect 10133 67222 12000 67224
rect 10133 67219 10199 67222
rect 11200 67192 12000 67222
rect 0 67146 800 67176
rect 1669 67146 1735 67149
rect 0 67144 1735 67146
rect 0 67088 1674 67144
rect 1730 67088 1735 67144
rect 0 67086 1735 67088
rect 0 67056 800 67086
rect 1669 67083 1735 67086
rect 2576 66944 2896 66945
rect 2576 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2576 66879 2896 66880
rect 5839 66944 6159 66945
rect 5839 66880 5847 66944
rect 5911 66880 5927 66944
rect 5991 66880 6007 66944
rect 6071 66880 6087 66944
rect 6151 66880 6159 66944
rect 5839 66879 6159 66880
rect 9103 66944 9423 66945
rect 9103 66880 9111 66944
rect 9175 66880 9191 66944
rect 9255 66880 9271 66944
rect 9335 66880 9351 66944
rect 9415 66880 9423 66944
rect 9103 66879 9423 66880
rect 0 66602 800 66632
rect 2773 66602 2839 66605
rect 0 66600 2839 66602
rect 0 66544 2778 66600
rect 2834 66544 2839 66600
rect 0 66542 2839 66544
rect 0 66512 800 66542
rect 2773 66539 2839 66542
rect 4207 66400 4527 66401
rect 4207 66336 4215 66400
rect 4279 66336 4295 66400
rect 4359 66336 4375 66400
rect 4439 66336 4455 66400
rect 4519 66336 4527 66400
rect 4207 66335 4527 66336
rect 7471 66400 7791 66401
rect 7471 66336 7479 66400
rect 7543 66336 7559 66400
rect 7623 66336 7639 66400
rect 7703 66336 7719 66400
rect 7783 66336 7791 66400
rect 7471 66335 7791 66336
rect 0 66194 800 66224
rect 1393 66194 1459 66197
rect 0 66192 1459 66194
rect 0 66136 1398 66192
rect 1454 66136 1459 66192
rect 0 66134 1459 66136
rect 0 66104 800 66134
rect 1393 66131 1459 66134
rect 10133 66058 10199 66061
rect 11200 66058 12000 66088
rect 10133 66056 12000 66058
rect 10133 66000 10138 66056
rect 10194 66000 12000 66056
rect 10133 65998 12000 66000
rect 10133 65995 10199 65998
rect 11200 65968 12000 65998
rect 2576 65856 2896 65857
rect 0 65786 800 65816
rect 2576 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2576 65791 2896 65792
rect 5839 65856 6159 65857
rect 5839 65792 5847 65856
rect 5911 65792 5927 65856
rect 5991 65792 6007 65856
rect 6071 65792 6087 65856
rect 6151 65792 6159 65856
rect 5839 65791 6159 65792
rect 9103 65856 9423 65857
rect 9103 65792 9111 65856
rect 9175 65792 9191 65856
rect 9255 65792 9271 65856
rect 9335 65792 9351 65856
rect 9415 65792 9423 65856
rect 9103 65791 9423 65792
rect 1945 65786 2011 65789
rect 0 65784 2011 65786
rect 0 65728 1950 65784
rect 2006 65728 2011 65784
rect 0 65726 2011 65728
rect 0 65696 800 65726
rect 1945 65723 2011 65726
rect 4207 65312 4527 65313
rect 0 65242 800 65272
rect 4207 65248 4215 65312
rect 4279 65248 4295 65312
rect 4359 65248 4375 65312
rect 4439 65248 4455 65312
rect 4519 65248 4527 65312
rect 4207 65247 4527 65248
rect 7471 65312 7791 65313
rect 7471 65248 7479 65312
rect 7543 65248 7559 65312
rect 7623 65248 7639 65312
rect 7703 65248 7719 65312
rect 7783 65248 7791 65312
rect 7471 65247 7791 65248
rect 1945 65242 2011 65245
rect 0 65240 2011 65242
rect 0 65184 1950 65240
rect 2006 65184 2011 65240
rect 0 65182 2011 65184
rect 0 65152 800 65182
rect 1945 65179 2011 65182
rect 10133 64970 10199 64973
rect 11200 64970 12000 65000
rect 10133 64968 12000 64970
rect 10133 64912 10138 64968
rect 10194 64912 12000 64968
rect 10133 64910 12000 64912
rect 10133 64907 10199 64910
rect 11200 64880 12000 64910
rect 0 64834 800 64864
rect 2313 64836 2379 64837
rect 0 64774 1456 64834
rect 0 64744 800 64774
rect 1396 64562 1456 64774
rect 2262 64772 2268 64836
rect 2332 64834 2379 64836
rect 2332 64832 2424 64834
rect 2374 64776 2424 64832
rect 2332 64774 2424 64776
rect 2332 64772 2379 64774
rect 2313 64771 2379 64772
rect 2576 64768 2896 64769
rect 2576 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2576 64703 2896 64704
rect 5839 64768 6159 64769
rect 5839 64704 5847 64768
rect 5911 64704 5927 64768
rect 5991 64704 6007 64768
rect 6071 64704 6087 64768
rect 6151 64704 6159 64768
rect 5839 64703 6159 64704
rect 9103 64768 9423 64769
rect 9103 64704 9111 64768
rect 9175 64704 9191 64768
rect 9255 64704 9271 64768
rect 9335 64704 9351 64768
rect 9415 64704 9423 64768
rect 9103 64703 9423 64704
rect 3141 64562 3207 64565
rect 1396 64560 3207 64562
rect 1396 64504 3146 64560
rect 3202 64504 3207 64560
rect 1396 64502 3207 64504
rect 3141 64499 3207 64502
rect 0 64426 800 64456
rect 3049 64426 3115 64429
rect 0 64424 3115 64426
rect 0 64368 3054 64424
rect 3110 64368 3115 64424
rect 0 64366 3115 64368
rect 0 64336 800 64366
rect 3049 64363 3115 64366
rect 4207 64224 4527 64225
rect 4207 64160 4215 64224
rect 4279 64160 4295 64224
rect 4359 64160 4375 64224
rect 4439 64160 4455 64224
rect 4519 64160 4527 64224
rect 4207 64159 4527 64160
rect 7471 64224 7791 64225
rect 7471 64160 7479 64224
rect 7543 64160 7559 64224
rect 7623 64160 7639 64224
rect 7703 64160 7719 64224
rect 7783 64160 7791 64224
rect 7471 64159 7791 64160
rect 0 64018 800 64048
rect 3969 64018 4035 64021
rect 0 64016 4035 64018
rect 0 63960 3974 64016
rect 4030 63960 4035 64016
rect 0 63958 4035 63960
rect 0 63928 800 63958
rect 3969 63955 4035 63958
rect 10133 63882 10199 63885
rect 11200 63882 12000 63912
rect 10133 63880 12000 63882
rect 10133 63824 10138 63880
rect 10194 63824 12000 63880
rect 10133 63822 12000 63824
rect 10133 63819 10199 63822
rect 11200 63792 12000 63822
rect 2576 63680 2896 63681
rect 2576 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2576 63615 2896 63616
rect 5839 63680 6159 63681
rect 5839 63616 5847 63680
rect 5911 63616 5927 63680
rect 5991 63616 6007 63680
rect 6071 63616 6087 63680
rect 6151 63616 6159 63680
rect 5839 63615 6159 63616
rect 9103 63680 9423 63681
rect 9103 63616 9111 63680
rect 9175 63616 9191 63680
rect 9255 63616 9271 63680
rect 9335 63616 9351 63680
rect 9415 63616 9423 63680
rect 9103 63615 9423 63616
rect 0 63474 800 63504
rect 1485 63474 1551 63477
rect 0 63472 1551 63474
rect 0 63416 1490 63472
rect 1546 63416 1551 63472
rect 0 63414 1551 63416
rect 0 63384 800 63414
rect 1485 63411 1551 63414
rect 4207 63136 4527 63137
rect 0 63066 800 63096
rect 4207 63072 4215 63136
rect 4279 63072 4295 63136
rect 4359 63072 4375 63136
rect 4439 63072 4455 63136
rect 4519 63072 4527 63136
rect 4207 63071 4527 63072
rect 7471 63136 7791 63137
rect 7471 63072 7479 63136
rect 7543 63072 7559 63136
rect 7623 63072 7639 63136
rect 7703 63072 7719 63136
rect 7783 63072 7791 63136
rect 7471 63071 7791 63072
rect 3969 63066 4035 63069
rect 0 63064 4035 63066
rect 0 63008 3974 63064
rect 4030 63008 4035 63064
rect 0 63006 4035 63008
rect 0 62976 800 63006
rect 3969 63003 4035 63006
rect 10133 62794 10199 62797
rect 11200 62794 12000 62824
rect 10133 62792 12000 62794
rect 10133 62736 10138 62792
rect 10194 62736 12000 62792
rect 10133 62734 12000 62736
rect 10133 62731 10199 62734
rect 11200 62704 12000 62734
rect 0 62658 800 62688
rect 1393 62658 1459 62661
rect 0 62656 1459 62658
rect 0 62600 1398 62656
rect 1454 62600 1459 62656
rect 0 62598 1459 62600
rect 0 62568 800 62598
rect 1393 62595 1459 62598
rect 2576 62592 2896 62593
rect 2576 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2576 62527 2896 62528
rect 5839 62592 6159 62593
rect 5839 62528 5847 62592
rect 5911 62528 5927 62592
rect 5991 62528 6007 62592
rect 6071 62528 6087 62592
rect 6151 62528 6159 62592
rect 5839 62527 6159 62528
rect 9103 62592 9423 62593
rect 9103 62528 9111 62592
rect 9175 62528 9191 62592
rect 9255 62528 9271 62592
rect 9335 62528 9351 62592
rect 9415 62528 9423 62592
rect 9103 62527 9423 62528
rect 0 62114 800 62144
rect 1485 62114 1551 62117
rect 0 62112 1551 62114
rect 0 62056 1490 62112
rect 1546 62056 1551 62112
rect 0 62054 1551 62056
rect 0 62024 800 62054
rect 1485 62051 1551 62054
rect 1945 62114 2011 62117
rect 2078 62114 2084 62116
rect 1945 62112 2084 62114
rect 1945 62056 1950 62112
rect 2006 62056 2084 62112
rect 1945 62054 2084 62056
rect 1945 62051 2011 62054
rect 2078 62052 2084 62054
rect 2148 62052 2154 62116
rect 4207 62048 4527 62049
rect 4207 61984 4215 62048
rect 4279 61984 4295 62048
rect 4359 61984 4375 62048
rect 4439 61984 4455 62048
rect 4519 61984 4527 62048
rect 4207 61983 4527 61984
rect 7471 62048 7791 62049
rect 7471 61984 7479 62048
rect 7543 61984 7559 62048
rect 7623 61984 7639 62048
rect 7703 61984 7719 62048
rect 7783 61984 7791 62048
rect 7471 61983 7791 61984
rect 0 61706 800 61736
rect 2221 61706 2287 61709
rect 0 61704 2287 61706
rect 0 61648 2226 61704
rect 2282 61648 2287 61704
rect 0 61646 2287 61648
rect 0 61616 800 61646
rect 2221 61643 2287 61646
rect 10133 61706 10199 61709
rect 11200 61706 12000 61736
rect 10133 61704 12000 61706
rect 10133 61648 10138 61704
rect 10194 61648 12000 61704
rect 10133 61646 12000 61648
rect 10133 61643 10199 61646
rect 11200 61616 12000 61646
rect 2262 61508 2268 61572
rect 2332 61570 2338 61572
rect 2405 61570 2471 61573
rect 2332 61568 2471 61570
rect 2332 61512 2410 61568
rect 2466 61512 2471 61568
rect 2332 61510 2471 61512
rect 2332 61508 2338 61510
rect 2405 61507 2471 61510
rect 2576 61504 2896 61505
rect 2576 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2576 61439 2896 61440
rect 5839 61504 6159 61505
rect 5839 61440 5847 61504
rect 5911 61440 5927 61504
rect 5991 61440 6007 61504
rect 6071 61440 6087 61504
rect 6151 61440 6159 61504
rect 5839 61439 6159 61440
rect 9103 61504 9423 61505
rect 9103 61440 9111 61504
rect 9175 61440 9191 61504
rect 9255 61440 9271 61504
rect 9335 61440 9351 61504
rect 9415 61440 9423 61504
rect 9103 61439 9423 61440
rect 0 61298 800 61328
rect 1393 61298 1459 61301
rect 0 61296 1459 61298
rect 0 61240 1398 61296
rect 1454 61240 1459 61296
rect 0 61238 1459 61240
rect 0 61208 800 61238
rect 1393 61235 1459 61238
rect 4207 60960 4527 60961
rect 4207 60896 4215 60960
rect 4279 60896 4295 60960
rect 4359 60896 4375 60960
rect 4439 60896 4455 60960
rect 4519 60896 4527 60960
rect 4207 60895 4527 60896
rect 7471 60960 7791 60961
rect 7471 60896 7479 60960
rect 7543 60896 7559 60960
rect 7623 60896 7639 60960
rect 7703 60896 7719 60960
rect 7783 60896 7791 60960
rect 7471 60895 7791 60896
rect 0 60754 800 60784
rect 1485 60754 1551 60757
rect 0 60752 1551 60754
rect 0 60696 1490 60752
rect 1546 60696 1551 60752
rect 0 60694 1551 60696
rect 0 60664 800 60694
rect 1485 60691 1551 60694
rect 10133 60618 10199 60621
rect 11200 60618 12000 60648
rect 10133 60616 12000 60618
rect 10133 60560 10138 60616
rect 10194 60560 12000 60616
rect 10133 60558 12000 60560
rect 10133 60555 10199 60558
rect 11200 60528 12000 60558
rect 2576 60416 2896 60417
rect 0 60346 800 60376
rect 2576 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2576 60351 2896 60352
rect 5839 60416 6159 60417
rect 5839 60352 5847 60416
rect 5911 60352 5927 60416
rect 5991 60352 6007 60416
rect 6071 60352 6087 60416
rect 6151 60352 6159 60416
rect 5839 60351 6159 60352
rect 9103 60416 9423 60417
rect 9103 60352 9111 60416
rect 9175 60352 9191 60416
rect 9255 60352 9271 60416
rect 9335 60352 9351 60416
rect 9415 60352 9423 60416
rect 9103 60351 9423 60352
rect 1393 60346 1459 60349
rect 0 60344 1459 60346
rect 0 60288 1398 60344
rect 1454 60288 1459 60344
rect 0 60286 1459 60288
rect 0 60256 800 60286
rect 1393 60283 1459 60286
rect 0 59938 800 59968
rect 1485 59938 1551 59941
rect 0 59936 1551 59938
rect 0 59880 1490 59936
rect 1546 59880 1551 59936
rect 0 59878 1551 59880
rect 0 59848 800 59878
rect 1485 59875 1551 59878
rect 4207 59872 4527 59873
rect 4207 59808 4215 59872
rect 4279 59808 4295 59872
rect 4359 59808 4375 59872
rect 4439 59808 4455 59872
rect 4519 59808 4527 59872
rect 4207 59807 4527 59808
rect 7471 59872 7791 59873
rect 7471 59808 7479 59872
rect 7543 59808 7559 59872
rect 7623 59808 7639 59872
rect 7703 59808 7719 59872
rect 7783 59808 7791 59872
rect 7471 59807 7791 59808
rect 0 59530 800 59560
rect 2221 59530 2287 59533
rect 0 59528 2287 59530
rect 0 59472 2226 59528
rect 2282 59472 2287 59528
rect 0 59470 2287 59472
rect 0 59440 800 59470
rect 2221 59467 2287 59470
rect 10133 59394 10199 59397
rect 11200 59394 12000 59424
rect 10133 59392 12000 59394
rect 10133 59336 10138 59392
rect 10194 59336 12000 59392
rect 10133 59334 12000 59336
rect 10133 59331 10199 59334
rect 2576 59328 2896 59329
rect 2576 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2576 59263 2896 59264
rect 5839 59328 6159 59329
rect 5839 59264 5847 59328
rect 5911 59264 5927 59328
rect 5991 59264 6007 59328
rect 6071 59264 6087 59328
rect 6151 59264 6159 59328
rect 5839 59263 6159 59264
rect 9103 59328 9423 59329
rect 9103 59264 9111 59328
rect 9175 59264 9191 59328
rect 9255 59264 9271 59328
rect 9335 59264 9351 59328
rect 9415 59264 9423 59328
rect 11200 59304 12000 59334
rect 9103 59263 9423 59264
rect 0 58986 800 59016
rect 1393 58986 1459 58989
rect 0 58984 1459 58986
rect 0 58928 1398 58984
rect 1454 58928 1459 58984
rect 0 58926 1459 58928
rect 0 58896 800 58926
rect 1393 58923 1459 58926
rect 4207 58784 4527 58785
rect 4207 58720 4215 58784
rect 4279 58720 4295 58784
rect 4359 58720 4375 58784
rect 4439 58720 4455 58784
rect 4519 58720 4527 58784
rect 4207 58719 4527 58720
rect 7471 58784 7791 58785
rect 7471 58720 7479 58784
rect 7543 58720 7559 58784
rect 7623 58720 7639 58784
rect 7703 58720 7719 58784
rect 7783 58720 7791 58784
rect 7471 58719 7791 58720
rect 0 58578 800 58608
rect 2773 58578 2839 58581
rect 0 58576 2839 58578
rect 0 58520 2778 58576
rect 2834 58520 2839 58576
rect 0 58518 2839 58520
rect 0 58488 800 58518
rect 2773 58515 2839 58518
rect 1669 58308 1735 58309
rect 1669 58306 1716 58308
rect 1624 58304 1716 58306
rect 1624 58248 1674 58304
rect 1624 58246 1716 58248
rect 1669 58244 1716 58246
rect 1780 58244 1786 58308
rect 10133 58306 10199 58309
rect 11200 58306 12000 58336
rect 10133 58304 12000 58306
rect 10133 58248 10138 58304
rect 10194 58248 12000 58304
rect 10133 58246 12000 58248
rect 1669 58243 1735 58244
rect 10133 58243 10199 58246
rect 2576 58240 2896 58241
rect 0 58170 800 58200
rect 2576 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2576 58175 2896 58176
rect 5839 58240 6159 58241
rect 5839 58176 5847 58240
rect 5911 58176 5927 58240
rect 5991 58176 6007 58240
rect 6071 58176 6087 58240
rect 6151 58176 6159 58240
rect 5839 58175 6159 58176
rect 9103 58240 9423 58241
rect 9103 58176 9111 58240
rect 9175 58176 9191 58240
rect 9255 58176 9271 58240
rect 9335 58176 9351 58240
rect 9415 58176 9423 58240
rect 11200 58216 12000 58246
rect 9103 58175 9423 58176
rect 1485 58170 1551 58173
rect 0 58168 1551 58170
rect 0 58112 1490 58168
rect 1546 58112 1551 58168
rect 0 58110 1551 58112
rect 0 58080 800 58110
rect 1485 58107 1551 58110
rect 4207 57696 4527 57697
rect 0 57626 800 57656
rect 4207 57632 4215 57696
rect 4279 57632 4295 57696
rect 4359 57632 4375 57696
rect 4439 57632 4455 57696
rect 4519 57632 4527 57696
rect 4207 57631 4527 57632
rect 7471 57696 7791 57697
rect 7471 57632 7479 57696
rect 7543 57632 7559 57696
rect 7623 57632 7639 57696
rect 7703 57632 7719 57696
rect 7783 57632 7791 57696
rect 7471 57631 7791 57632
rect 2497 57626 2563 57629
rect 0 57624 2563 57626
rect 0 57568 2502 57624
rect 2558 57568 2563 57624
rect 0 57566 2563 57568
rect 0 57536 800 57566
rect 2497 57563 2563 57566
rect 3141 57354 3207 57357
rect 1350 57352 3207 57354
rect 1350 57296 3146 57352
rect 3202 57296 3207 57352
rect 1350 57294 3207 57296
rect 0 57218 800 57248
rect 1350 57218 1410 57294
rect 3141 57291 3207 57294
rect 0 57158 1410 57218
rect 10133 57218 10199 57221
rect 11200 57218 12000 57248
rect 10133 57216 12000 57218
rect 10133 57160 10138 57216
rect 10194 57160 12000 57216
rect 10133 57158 12000 57160
rect 0 57128 800 57158
rect 10133 57155 10199 57158
rect 2576 57152 2896 57153
rect 2576 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2576 57087 2896 57088
rect 5839 57152 6159 57153
rect 5839 57088 5847 57152
rect 5911 57088 5927 57152
rect 5991 57088 6007 57152
rect 6071 57088 6087 57152
rect 6151 57088 6159 57152
rect 5839 57087 6159 57088
rect 9103 57152 9423 57153
rect 9103 57088 9111 57152
rect 9175 57088 9191 57152
rect 9255 57088 9271 57152
rect 9335 57088 9351 57152
rect 9415 57088 9423 57152
rect 11200 57128 12000 57158
rect 9103 57087 9423 57088
rect 0 56810 800 56840
rect 2497 56810 2563 56813
rect 0 56808 2563 56810
rect 0 56752 2502 56808
rect 2558 56752 2563 56808
rect 0 56750 2563 56752
rect 0 56720 800 56750
rect 2497 56747 2563 56750
rect 3049 56676 3115 56677
rect 2998 56674 3004 56676
rect 2958 56614 3004 56674
rect 3068 56672 3115 56676
rect 3110 56616 3115 56672
rect 2998 56612 3004 56614
rect 3068 56612 3115 56616
rect 3049 56611 3115 56612
rect 4207 56608 4527 56609
rect 4207 56544 4215 56608
rect 4279 56544 4295 56608
rect 4359 56544 4375 56608
rect 4439 56544 4455 56608
rect 4519 56544 4527 56608
rect 4207 56543 4527 56544
rect 7471 56608 7791 56609
rect 7471 56544 7479 56608
rect 7543 56544 7559 56608
rect 7623 56544 7639 56608
rect 7703 56544 7719 56608
rect 7783 56544 7791 56608
rect 7471 56543 7791 56544
rect 0 56266 800 56296
rect 2313 56266 2379 56269
rect 0 56264 2379 56266
rect 0 56208 2318 56264
rect 2374 56208 2379 56264
rect 0 56206 2379 56208
rect 0 56176 800 56206
rect 2313 56203 2379 56206
rect 4654 56204 4660 56268
rect 4724 56266 4730 56268
rect 4797 56266 4863 56269
rect 4724 56264 4863 56266
rect 4724 56208 4802 56264
rect 4858 56208 4863 56264
rect 4724 56206 4863 56208
rect 4724 56204 4730 56206
rect 4797 56203 4863 56206
rect 10133 56130 10199 56133
rect 11200 56130 12000 56160
rect 10133 56128 12000 56130
rect 10133 56072 10138 56128
rect 10194 56072 12000 56128
rect 10133 56070 12000 56072
rect 10133 56067 10199 56070
rect 2576 56064 2896 56065
rect 2576 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2576 55999 2896 56000
rect 5839 56064 6159 56065
rect 5839 56000 5847 56064
rect 5911 56000 5927 56064
rect 5991 56000 6007 56064
rect 6071 56000 6087 56064
rect 6151 56000 6159 56064
rect 5839 55999 6159 56000
rect 9103 56064 9423 56065
rect 9103 56000 9111 56064
rect 9175 56000 9191 56064
rect 9255 56000 9271 56064
rect 9335 56000 9351 56064
rect 9415 56000 9423 56064
rect 11200 56040 12000 56070
rect 9103 55999 9423 56000
rect 0 55858 800 55888
rect 1485 55858 1551 55861
rect 0 55856 1551 55858
rect 0 55800 1490 55856
rect 1546 55800 1551 55856
rect 0 55798 1551 55800
rect 0 55768 800 55798
rect 1485 55795 1551 55798
rect 3182 55796 3188 55860
rect 3252 55858 3258 55860
rect 3601 55858 3667 55861
rect 3252 55856 3667 55858
rect 3252 55800 3606 55856
rect 3662 55800 3667 55856
rect 3252 55798 3667 55800
rect 3252 55796 3258 55798
rect 3601 55795 3667 55798
rect 4207 55520 4527 55521
rect 0 55450 800 55480
rect 4207 55456 4215 55520
rect 4279 55456 4295 55520
rect 4359 55456 4375 55520
rect 4439 55456 4455 55520
rect 4519 55456 4527 55520
rect 4207 55455 4527 55456
rect 7471 55520 7791 55521
rect 7471 55456 7479 55520
rect 7543 55456 7559 55520
rect 7623 55456 7639 55520
rect 7703 55456 7719 55520
rect 7783 55456 7791 55520
rect 7471 55455 7791 55456
rect 1485 55450 1551 55453
rect 0 55448 1551 55450
rect 0 55392 1490 55448
rect 1546 55392 1551 55448
rect 0 55390 1551 55392
rect 0 55360 800 55390
rect 1485 55387 1551 55390
rect 1158 55252 1164 55316
rect 1228 55314 1234 55316
rect 1393 55314 1459 55317
rect 1228 55312 1459 55314
rect 1228 55256 1398 55312
rect 1454 55256 1459 55312
rect 1228 55254 1459 55256
rect 1228 55252 1234 55254
rect 1393 55251 1459 55254
rect 0 55042 800 55072
rect 2221 55042 2287 55045
rect 0 55040 2287 55042
rect 0 54984 2226 55040
rect 2282 54984 2287 55040
rect 0 54982 2287 54984
rect 0 54952 800 54982
rect 2221 54979 2287 54982
rect 10133 55042 10199 55045
rect 11200 55042 12000 55072
rect 10133 55040 12000 55042
rect 10133 54984 10138 55040
rect 10194 54984 12000 55040
rect 10133 54982 12000 54984
rect 10133 54979 10199 54982
rect 2576 54976 2896 54977
rect 2576 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2576 54911 2896 54912
rect 5839 54976 6159 54977
rect 5839 54912 5847 54976
rect 5911 54912 5927 54976
rect 5991 54912 6007 54976
rect 6071 54912 6087 54976
rect 6151 54912 6159 54976
rect 5839 54911 6159 54912
rect 9103 54976 9423 54977
rect 9103 54912 9111 54976
rect 9175 54912 9191 54976
rect 9255 54912 9271 54976
rect 9335 54912 9351 54976
rect 9415 54912 9423 54976
rect 11200 54952 12000 54982
rect 9103 54911 9423 54912
rect 3366 54708 3372 54772
rect 3436 54770 3442 54772
rect 3969 54770 4035 54773
rect 3436 54768 4035 54770
rect 3436 54712 3974 54768
rect 4030 54712 4035 54768
rect 3436 54710 4035 54712
rect 3436 54708 3442 54710
rect 3969 54707 4035 54710
rect 0 54498 800 54528
rect 1485 54498 1551 54501
rect 0 54496 1551 54498
rect 0 54440 1490 54496
rect 1546 54440 1551 54496
rect 0 54438 1551 54440
rect 0 54408 800 54438
rect 1485 54435 1551 54438
rect 4207 54432 4527 54433
rect 4207 54368 4215 54432
rect 4279 54368 4295 54432
rect 4359 54368 4375 54432
rect 4439 54368 4455 54432
rect 4519 54368 4527 54432
rect 4207 54367 4527 54368
rect 7471 54432 7791 54433
rect 7471 54368 7479 54432
rect 7543 54368 7559 54432
rect 7623 54368 7639 54432
rect 7703 54368 7719 54432
rect 7783 54368 7791 54432
rect 7471 54367 7791 54368
rect 0 54090 800 54120
rect 2221 54090 2287 54093
rect 0 54088 2287 54090
rect 0 54032 2226 54088
rect 2282 54032 2287 54088
rect 0 54030 2287 54032
rect 0 54000 800 54030
rect 2221 54027 2287 54030
rect 2037 53954 2103 53957
rect 10133 53954 10199 53957
rect 11200 53954 12000 53984
rect 2037 53952 2146 53954
rect 2037 53896 2042 53952
rect 2098 53896 2146 53952
rect 2037 53891 2146 53896
rect 10133 53952 12000 53954
rect 10133 53896 10138 53952
rect 10194 53896 12000 53952
rect 10133 53894 12000 53896
rect 10133 53891 10199 53894
rect 0 53682 800 53712
rect 1393 53682 1459 53685
rect 0 53680 1459 53682
rect 0 53624 1398 53680
rect 1454 53624 1459 53680
rect 0 53622 1459 53624
rect 2086 53682 2146 53891
rect 2576 53888 2896 53889
rect 2576 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2576 53823 2896 53824
rect 5839 53888 6159 53889
rect 5839 53824 5847 53888
rect 5911 53824 5927 53888
rect 5991 53824 6007 53888
rect 6071 53824 6087 53888
rect 6151 53824 6159 53888
rect 5839 53823 6159 53824
rect 9103 53888 9423 53889
rect 9103 53824 9111 53888
rect 9175 53824 9191 53888
rect 9255 53824 9271 53888
rect 9335 53824 9351 53888
rect 9415 53824 9423 53888
rect 11200 53864 12000 53894
rect 9103 53823 9423 53824
rect 2221 53682 2287 53685
rect 5441 53684 5507 53685
rect 2086 53680 2287 53682
rect 2086 53624 2226 53680
rect 2282 53624 2287 53680
rect 2086 53622 2287 53624
rect 0 53592 800 53622
rect 1393 53619 1459 53622
rect 2221 53619 2287 53622
rect 5390 53620 5396 53684
rect 5460 53682 5507 53684
rect 5460 53680 5552 53682
rect 5502 53624 5552 53680
rect 5460 53622 5552 53624
rect 5460 53620 5507 53622
rect 5441 53619 5507 53620
rect 1945 53410 2011 53413
rect 2262 53410 2268 53412
rect 1945 53408 2268 53410
rect 1945 53352 1950 53408
rect 2006 53352 2268 53408
rect 1945 53350 2268 53352
rect 1945 53347 2011 53350
rect 2262 53348 2268 53350
rect 2332 53348 2338 53412
rect 4207 53344 4527 53345
rect 4207 53280 4215 53344
rect 4279 53280 4295 53344
rect 4359 53280 4375 53344
rect 4439 53280 4455 53344
rect 4519 53280 4527 53344
rect 4207 53279 4527 53280
rect 7471 53344 7791 53345
rect 7471 53280 7479 53344
rect 7543 53280 7559 53344
rect 7623 53280 7639 53344
rect 7703 53280 7719 53344
rect 7783 53280 7791 53344
rect 7471 53279 7791 53280
rect 0 53138 800 53168
rect 2313 53138 2379 53141
rect 0 53136 2379 53138
rect 0 53080 2318 53136
rect 2374 53080 2379 53136
rect 0 53078 2379 53080
rect 0 53048 800 53078
rect 2313 53075 2379 53078
rect 4838 53076 4844 53140
rect 4908 53138 4914 53140
rect 5349 53138 5415 53141
rect 4908 53136 5415 53138
rect 4908 53080 5354 53136
rect 5410 53080 5415 53136
rect 4908 53078 5415 53080
rect 4908 53076 4914 53078
rect 5349 53075 5415 53078
rect 2576 52800 2896 52801
rect 0 52730 800 52760
rect 2576 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2576 52735 2896 52736
rect 5839 52800 6159 52801
rect 5839 52736 5847 52800
rect 5911 52736 5927 52800
rect 5991 52736 6007 52800
rect 6071 52736 6087 52800
rect 6151 52736 6159 52800
rect 5839 52735 6159 52736
rect 9103 52800 9423 52801
rect 9103 52736 9111 52800
rect 9175 52736 9191 52800
rect 9255 52736 9271 52800
rect 9335 52736 9351 52800
rect 9415 52736 9423 52800
rect 9103 52735 9423 52736
rect 1485 52730 1551 52733
rect 0 52728 1551 52730
rect 0 52672 1490 52728
rect 1546 52672 1551 52728
rect 0 52670 1551 52672
rect 0 52640 800 52670
rect 1485 52667 1551 52670
rect 10133 52730 10199 52733
rect 11200 52730 12000 52760
rect 10133 52728 12000 52730
rect 10133 52672 10138 52728
rect 10194 52672 12000 52728
rect 10133 52670 12000 52672
rect 10133 52667 10199 52670
rect 11200 52640 12000 52670
rect 0 52322 800 52352
rect 2957 52322 3023 52325
rect 0 52320 3023 52322
rect 0 52264 2962 52320
rect 3018 52264 3023 52320
rect 0 52262 3023 52264
rect 0 52232 800 52262
rect 2957 52259 3023 52262
rect 4207 52256 4527 52257
rect 4207 52192 4215 52256
rect 4279 52192 4295 52256
rect 4359 52192 4375 52256
rect 4439 52192 4455 52256
rect 4519 52192 4527 52256
rect 4207 52191 4527 52192
rect 7471 52256 7791 52257
rect 7471 52192 7479 52256
rect 7543 52192 7559 52256
rect 7623 52192 7639 52256
rect 7703 52192 7719 52256
rect 7783 52192 7791 52256
rect 7471 52191 7791 52192
rect 0 51778 800 51808
rect 1393 51778 1459 51781
rect 0 51776 1459 51778
rect 0 51720 1398 51776
rect 1454 51720 1459 51776
rect 0 51718 1459 51720
rect 0 51688 800 51718
rect 1393 51715 1459 51718
rect 2576 51712 2896 51713
rect 2576 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2576 51647 2896 51648
rect 5839 51712 6159 51713
rect 5839 51648 5847 51712
rect 5911 51648 5927 51712
rect 5991 51648 6007 51712
rect 6071 51648 6087 51712
rect 6151 51648 6159 51712
rect 5839 51647 6159 51648
rect 9103 51712 9423 51713
rect 9103 51648 9111 51712
rect 9175 51648 9191 51712
rect 9255 51648 9271 51712
rect 9335 51648 9351 51712
rect 9415 51648 9423 51712
rect 9103 51647 9423 51648
rect 4797 51644 4863 51645
rect 4797 51642 4844 51644
rect 4752 51640 4844 51642
rect 4752 51584 4802 51640
rect 4752 51582 4844 51584
rect 4797 51580 4844 51582
rect 4908 51580 4914 51644
rect 10133 51642 10199 51645
rect 11200 51642 12000 51672
rect 10133 51640 12000 51642
rect 10133 51584 10138 51640
rect 10194 51584 12000 51640
rect 10133 51582 12000 51584
rect 4797 51579 4863 51580
rect 10133 51579 10199 51582
rect 11200 51552 12000 51582
rect 1577 51506 1643 51509
rect 3785 51506 3851 51509
rect 1577 51504 3851 51506
rect 1577 51448 1582 51504
rect 1638 51448 3790 51504
rect 3846 51448 3851 51504
rect 1577 51446 3851 51448
rect 1577 51443 1643 51446
rect 3785 51443 3851 51446
rect 0 51370 800 51400
rect 1485 51370 1551 51373
rect 2129 51370 2195 51373
rect 5349 51370 5415 51373
rect 0 51368 1551 51370
rect 0 51312 1490 51368
rect 1546 51312 1551 51368
rect 0 51310 1551 51312
rect 0 51280 800 51310
rect 1485 51307 1551 51310
rect 2086 51368 2195 51370
rect 2086 51312 2134 51368
rect 2190 51312 2195 51368
rect 2086 51307 2195 51312
rect 5214 51368 5415 51370
rect 5214 51312 5354 51368
rect 5410 51312 5415 51368
rect 5214 51310 5415 51312
rect 1301 51234 1367 51237
rect 1301 51232 1594 51234
rect 1301 51176 1306 51232
rect 1362 51176 1594 51232
rect 1301 51174 1594 51176
rect 1301 51171 1367 51174
rect 1534 51101 1594 51174
rect 1534 51096 1643 51101
rect 1534 51040 1582 51096
rect 1638 51040 1643 51096
rect 1534 51038 1643 51040
rect 1577 51035 1643 51038
rect 1945 51098 2011 51101
rect 2086 51098 2146 51307
rect 2313 51236 2379 51237
rect 2262 51172 2268 51236
rect 2332 51234 2379 51236
rect 4981 51234 5047 51237
rect 2332 51232 2424 51234
rect 2374 51176 2424 51232
rect 2332 51174 2424 51176
rect 4846 51232 5047 51234
rect 4846 51176 4986 51232
rect 5042 51176 5047 51232
rect 4846 51174 5047 51176
rect 2332 51172 2379 51174
rect 2313 51171 2379 51172
rect 4207 51168 4527 51169
rect 4207 51104 4215 51168
rect 4279 51104 4295 51168
rect 4359 51104 4375 51168
rect 4439 51104 4455 51168
rect 4519 51104 4527 51168
rect 4207 51103 4527 51104
rect 1945 51096 2146 51098
rect 1945 51040 1950 51096
rect 2006 51040 2146 51096
rect 3969 51090 4035 51093
rect 1945 51038 2146 51040
rect 3926 51088 4035 51090
rect 1945 51035 2011 51038
rect 3926 51032 3974 51088
rect 4030 51032 4035 51088
rect 3926 51027 4035 51032
rect 0 50962 800 50992
rect 3926 50962 3986 51027
rect 0 50902 3986 50962
rect 4846 50965 4906 51174
rect 4981 51171 5047 51174
rect 4846 50960 4955 50965
rect 4846 50904 4894 50960
rect 4950 50904 4955 50960
rect 4846 50902 4955 50904
rect 5214 50962 5274 51310
rect 5349 51307 5415 51310
rect 7471 51168 7791 51169
rect 7471 51104 7479 51168
rect 7543 51104 7559 51168
rect 7623 51104 7639 51168
rect 7703 51104 7719 51168
rect 7783 51104 7791 51168
rect 7471 51103 7791 51104
rect 5441 51100 5507 51101
rect 5390 51036 5396 51100
rect 5460 51098 5507 51100
rect 5460 51096 5552 51098
rect 5502 51040 5552 51096
rect 5460 51038 5552 51040
rect 5460 51036 5507 51038
rect 5441 51035 5507 51036
rect 5349 50962 5415 50965
rect 5214 50960 5415 50962
rect 5214 50904 5354 50960
rect 5410 50904 5415 50960
rect 5214 50902 5415 50904
rect 0 50872 800 50902
rect 4889 50899 4955 50902
rect 5349 50899 5415 50902
rect 2957 50826 3023 50829
rect 3233 50826 3299 50829
rect 3601 50826 3667 50829
rect 2957 50824 3299 50826
rect 2957 50768 2962 50824
rect 3018 50768 3238 50824
rect 3294 50768 3299 50824
rect 2957 50766 3299 50768
rect 2957 50763 3023 50766
rect 3233 50763 3299 50766
rect 3558 50824 3667 50826
rect 3558 50768 3606 50824
rect 3662 50768 3667 50824
rect 3558 50763 3667 50768
rect 3049 50690 3115 50693
rect 3182 50690 3188 50692
rect 3049 50688 3188 50690
rect 3049 50632 3054 50688
rect 3110 50632 3188 50688
rect 3049 50630 3188 50632
rect 3049 50627 3115 50630
rect 3182 50628 3188 50630
rect 3252 50628 3258 50692
rect 2576 50624 2896 50625
rect 2576 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2576 50559 2896 50560
rect 0 50418 800 50448
rect 3417 50418 3483 50421
rect 0 50416 3483 50418
rect 0 50360 3422 50416
rect 3478 50360 3483 50416
rect 0 50358 3483 50360
rect 0 50328 800 50358
rect 3417 50355 3483 50358
rect 1761 50282 1827 50285
rect 2497 50282 2563 50285
rect 1761 50280 2563 50282
rect 1761 50224 1766 50280
rect 1822 50224 2502 50280
rect 2558 50224 2563 50280
rect 1761 50222 2563 50224
rect 1761 50219 1827 50222
rect 2497 50219 2563 50222
rect 3325 50282 3391 50285
rect 3558 50282 3618 50763
rect 5839 50624 6159 50625
rect 5839 50560 5847 50624
rect 5911 50560 5927 50624
rect 5991 50560 6007 50624
rect 6071 50560 6087 50624
rect 6151 50560 6159 50624
rect 5839 50559 6159 50560
rect 9103 50624 9423 50625
rect 9103 50560 9111 50624
rect 9175 50560 9191 50624
rect 9255 50560 9271 50624
rect 9335 50560 9351 50624
rect 9415 50560 9423 50624
rect 9103 50559 9423 50560
rect 10133 50554 10199 50557
rect 11200 50554 12000 50584
rect 10133 50552 12000 50554
rect 10133 50496 10138 50552
rect 10194 50496 12000 50552
rect 10133 50494 12000 50496
rect 10133 50491 10199 50494
rect 11200 50464 12000 50494
rect 3325 50280 3618 50282
rect 3325 50224 3330 50280
rect 3386 50224 3618 50280
rect 3325 50222 3618 50224
rect 3325 50219 3391 50222
rect 4207 50080 4527 50081
rect 0 50010 800 50040
rect 4207 50016 4215 50080
rect 4279 50016 4295 50080
rect 4359 50016 4375 50080
rect 4439 50016 4455 50080
rect 4519 50016 4527 50080
rect 4207 50015 4527 50016
rect 7471 50080 7791 50081
rect 7471 50016 7479 50080
rect 7543 50016 7559 50080
rect 7623 50016 7639 50080
rect 7703 50016 7719 50080
rect 7783 50016 7791 50080
rect 7471 50015 7791 50016
rect 2497 50010 2563 50013
rect 0 50008 2563 50010
rect 0 49952 2502 50008
rect 2558 49952 2563 50008
rect 0 49950 2563 49952
rect 0 49920 800 49950
rect 2497 49947 2563 49950
rect 0 49602 800 49632
rect 2221 49602 2287 49605
rect 0 49600 2287 49602
rect 0 49544 2226 49600
rect 2282 49544 2287 49600
rect 0 49542 2287 49544
rect 0 49512 800 49542
rect 2221 49539 2287 49542
rect 2576 49536 2896 49537
rect 2576 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2576 49471 2896 49472
rect 5839 49536 6159 49537
rect 5839 49472 5847 49536
rect 5911 49472 5927 49536
rect 5991 49472 6007 49536
rect 6071 49472 6087 49536
rect 6151 49472 6159 49536
rect 5839 49471 6159 49472
rect 9103 49536 9423 49537
rect 9103 49472 9111 49536
rect 9175 49472 9191 49536
rect 9255 49472 9271 49536
rect 9335 49472 9351 49536
rect 9415 49472 9423 49536
rect 9103 49471 9423 49472
rect 10133 49466 10199 49469
rect 11200 49466 12000 49496
rect 10133 49464 12000 49466
rect 10133 49408 10138 49464
rect 10194 49408 12000 49464
rect 10133 49406 12000 49408
rect 10133 49403 10199 49406
rect 11200 49376 12000 49406
rect 3233 49330 3299 49333
rect 3366 49330 3372 49332
rect 3233 49328 3372 49330
rect 3233 49272 3238 49328
rect 3294 49272 3372 49328
rect 3233 49270 3372 49272
rect 3233 49267 3299 49270
rect 3366 49268 3372 49270
rect 3436 49268 3442 49332
rect 0 49194 800 49224
rect 1485 49194 1551 49197
rect 0 49192 1551 49194
rect 0 49136 1490 49192
rect 1546 49136 1551 49192
rect 0 49134 1551 49136
rect 0 49104 800 49134
rect 1485 49131 1551 49134
rect 4207 48992 4527 48993
rect 4207 48928 4215 48992
rect 4279 48928 4295 48992
rect 4359 48928 4375 48992
rect 4439 48928 4455 48992
rect 4519 48928 4527 48992
rect 4207 48927 4527 48928
rect 7471 48992 7791 48993
rect 7471 48928 7479 48992
rect 7543 48928 7559 48992
rect 7623 48928 7639 48992
rect 7703 48928 7719 48992
rect 7783 48928 7791 48992
rect 7471 48927 7791 48928
rect 4429 48786 4495 48789
rect 4654 48786 4660 48788
rect 4429 48784 4660 48786
rect 4429 48728 4434 48784
rect 4490 48728 4660 48784
rect 4429 48726 4660 48728
rect 4429 48723 4495 48726
rect 4654 48724 4660 48726
rect 4724 48724 4730 48788
rect 6678 48724 6684 48788
rect 6748 48786 6754 48788
rect 6821 48786 6887 48789
rect 6748 48784 6887 48786
rect 6748 48728 6826 48784
rect 6882 48728 6887 48784
rect 6748 48726 6887 48728
rect 6748 48724 6754 48726
rect 6821 48723 6887 48726
rect 0 48650 800 48680
rect 2221 48650 2287 48653
rect 0 48648 2287 48650
rect 0 48592 2226 48648
rect 2282 48592 2287 48648
rect 0 48590 2287 48592
rect 0 48560 800 48590
rect 2221 48587 2287 48590
rect 2576 48448 2896 48449
rect 2576 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2576 48383 2896 48384
rect 5839 48448 6159 48449
rect 5839 48384 5847 48448
rect 5911 48384 5927 48448
rect 5991 48384 6007 48448
rect 6071 48384 6087 48448
rect 6151 48384 6159 48448
rect 5839 48383 6159 48384
rect 9103 48448 9423 48449
rect 9103 48384 9111 48448
rect 9175 48384 9191 48448
rect 9255 48384 9271 48448
rect 9335 48384 9351 48448
rect 9415 48384 9423 48448
rect 9103 48383 9423 48384
rect 10133 48378 10199 48381
rect 11200 48378 12000 48408
rect 10133 48376 12000 48378
rect 10133 48320 10138 48376
rect 10194 48320 12000 48376
rect 10133 48318 12000 48320
rect 10133 48315 10199 48318
rect 11200 48288 12000 48318
rect 0 48242 800 48272
rect 1485 48242 1551 48245
rect 0 48240 1551 48242
rect 0 48184 1490 48240
rect 1546 48184 1551 48240
rect 0 48182 1551 48184
rect 0 48152 800 48182
rect 1485 48179 1551 48182
rect 3734 48180 3740 48244
rect 3804 48242 3810 48244
rect 4429 48242 4495 48245
rect 3804 48240 4495 48242
rect 3804 48184 4434 48240
rect 4490 48184 4495 48240
rect 3804 48182 4495 48184
rect 3804 48180 3810 48182
rect 4429 48179 4495 48182
rect 4521 48106 4587 48109
rect 4654 48106 4660 48108
rect 4521 48104 4660 48106
rect 4521 48048 4526 48104
rect 4582 48048 4660 48104
rect 4521 48046 4660 48048
rect 4521 48043 4587 48046
rect 4654 48044 4660 48046
rect 4724 48044 4730 48108
rect 4207 47904 4527 47905
rect 0 47834 800 47864
rect 4207 47840 4215 47904
rect 4279 47840 4295 47904
rect 4359 47840 4375 47904
rect 4439 47840 4455 47904
rect 4519 47840 4527 47904
rect 4207 47839 4527 47840
rect 7471 47904 7791 47905
rect 7471 47840 7479 47904
rect 7543 47840 7559 47904
rect 7623 47840 7639 47904
rect 7703 47840 7719 47904
rect 7783 47840 7791 47904
rect 7471 47839 7791 47840
rect 1485 47834 1551 47837
rect 0 47832 1551 47834
rect 0 47776 1490 47832
rect 1546 47776 1551 47832
rect 0 47774 1551 47776
rect 0 47744 800 47774
rect 1485 47771 1551 47774
rect 2865 47698 2931 47701
rect 3877 47698 3943 47701
rect 2865 47696 3943 47698
rect 2865 47640 2870 47696
rect 2926 47640 3882 47696
rect 3938 47640 3943 47696
rect 2865 47638 3943 47640
rect 2865 47635 2931 47638
rect 3877 47635 3943 47638
rect 2576 47360 2896 47361
rect 0 47290 800 47320
rect 2576 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2576 47295 2896 47296
rect 5839 47360 6159 47361
rect 5839 47296 5847 47360
rect 5911 47296 5927 47360
rect 5991 47296 6007 47360
rect 6071 47296 6087 47360
rect 6151 47296 6159 47360
rect 5839 47295 6159 47296
rect 9103 47360 9423 47361
rect 9103 47296 9111 47360
rect 9175 47296 9191 47360
rect 9255 47296 9271 47360
rect 9335 47296 9351 47360
rect 9415 47296 9423 47360
rect 9103 47295 9423 47296
rect 2221 47290 2287 47293
rect 0 47288 2287 47290
rect 0 47232 2226 47288
rect 2282 47232 2287 47288
rect 0 47230 2287 47232
rect 0 47200 800 47230
rect 2221 47227 2287 47230
rect 10133 47290 10199 47293
rect 11200 47290 12000 47320
rect 10133 47288 12000 47290
rect 10133 47232 10138 47288
rect 10194 47232 12000 47288
rect 10133 47230 12000 47232
rect 10133 47227 10199 47230
rect 11200 47200 12000 47230
rect 0 46882 800 46912
rect 1485 46882 1551 46885
rect 0 46880 1551 46882
rect 0 46824 1490 46880
rect 1546 46824 1551 46880
rect 0 46822 1551 46824
rect 0 46792 800 46822
rect 1485 46819 1551 46822
rect 2497 46882 2563 46885
rect 2998 46882 3004 46884
rect 2497 46880 3004 46882
rect 2497 46824 2502 46880
rect 2558 46824 3004 46880
rect 2497 46822 3004 46824
rect 2497 46819 2563 46822
rect 2998 46820 3004 46822
rect 3068 46820 3074 46884
rect 4207 46816 4527 46817
rect 4207 46752 4215 46816
rect 4279 46752 4295 46816
rect 4359 46752 4375 46816
rect 4439 46752 4455 46816
rect 4519 46752 4527 46816
rect 4207 46751 4527 46752
rect 7471 46816 7791 46817
rect 7471 46752 7479 46816
rect 7543 46752 7559 46816
rect 7623 46752 7639 46816
rect 7703 46752 7719 46816
rect 7783 46752 7791 46816
rect 7471 46751 7791 46752
rect 0 46474 800 46504
rect 3049 46474 3115 46477
rect 0 46472 3115 46474
rect 0 46416 3054 46472
rect 3110 46416 3115 46472
rect 0 46414 3115 46416
rect 0 46384 800 46414
rect 3049 46411 3115 46414
rect 6729 46340 6795 46341
rect 6678 46276 6684 46340
rect 6748 46338 6795 46340
rect 6748 46336 6840 46338
rect 6790 46280 6840 46336
rect 6748 46278 6840 46280
rect 6748 46276 6795 46278
rect 6729 46275 6795 46276
rect 2576 46272 2896 46273
rect 2576 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2576 46207 2896 46208
rect 5839 46272 6159 46273
rect 5839 46208 5847 46272
rect 5911 46208 5927 46272
rect 5991 46208 6007 46272
rect 6071 46208 6087 46272
rect 6151 46208 6159 46272
rect 5839 46207 6159 46208
rect 9103 46272 9423 46273
rect 9103 46208 9111 46272
rect 9175 46208 9191 46272
rect 9255 46208 9271 46272
rect 9335 46208 9351 46272
rect 9415 46208 9423 46272
rect 9103 46207 9423 46208
rect 1485 46066 1551 46069
rect 2262 46066 2268 46068
rect 1485 46064 2268 46066
rect 1485 46008 1490 46064
rect 1546 46008 2268 46064
rect 1485 46006 2268 46008
rect 1485 46003 1551 46006
rect 2262 46004 2268 46006
rect 2332 46004 2338 46068
rect 10133 46066 10199 46069
rect 11200 46066 12000 46096
rect 10133 46064 12000 46066
rect 10133 46008 10138 46064
rect 10194 46008 12000 46064
rect 10133 46006 12000 46008
rect 10133 46003 10199 46006
rect 11200 45976 12000 46006
rect 0 45930 800 45960
rect 2221 45930 2287 45933
rect 0 45928 2287 45930
rect 0 45872 2226 45928
rect 2282 45872 2287 45928
rect 0 45870 2287 45872
rect 0 45840 800 45870
rect 2221 45867 2287 45870
rect 4207 45728 4527 45729
rect 4207 45664 4215 45728
rect 4279 45664 4295 45728
rect 4359 45664 4375 45728
rect 4439 45664 4455 45728
rect 4519 45664 4527 45728
rect 4207 45663 4527 45664
rect 7471 45728 7791 45729
rect 7471 45664 7479 45728
rect 7543 45664 7559 45728
rect 7623 45664 7639 45728
rect 7703 45664 7719 45728
rect 7783 45664 7791 45728
rect 7471 45663 7791 45664
rect 0 45522 800 45552
rect 1301 45522 1367 45525
rect 0 45520 1367 45522
rect 0 45464 1306 45520
rect 1362 45464 1367 45520
rect 0 45462 1367 45464
rect 0 45432 800 45462
rect 1301 45459 1367 45462
rect 2576 45184 2896 45185
rect 0 45114 800 45144
rect 2576 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2576 45119 2896 45120
rect 5839 45184 6159 45185
rect 5839 45120 5847 45184
rect 5911 45120 5927 45184
rect 5991 45120 6007 45184
rect 6071 45120 6087 45184
rect 6151 45120 6159 45184
rect 5839 45119 6159 45120
rect 9103 45184 9423 45185
rect 9103 45120 9111 45184
rect 9175 45120 9191 45184
rect 9255 45120 9271 45184
rect 9335 45120 9351 45184
rect 9415 45120 9423 45184
rect 9103 45119 9423 45120
rect 1393 45114 1459 45117
rect 0 45112 1459 45114
rect 0 45056 1398 45112
rect 1454 45056 1459 45112
rect 0 45054 1459 45056
rect 0 45024 800 45054
rect 1393 45051 1459 45054
rect 10133 44978 10199 44981
rect 11200 44978 12000 45008
rect 10133 44976 12000 44978
rect 10133 44920 10138 44976
rect 10194 44920 12000 44976
rect 10133 44918 12000 44920
rect 10133 44915 10199 44918
rect 11200 44888 12000 44918
rect 1577 44842 1643 44845
rect 2221 44842 2287 44845
rect 1577 44840 2287 44842
rect 1577 44784 1582 44840
rect 1638 44784 2226 44840
rect 2282 44784 2287 44840
rect 1577 44782 2287 44784
rect 1577 44779 1643 44782
rect 2221 44779 2287 44782
rect 0 44706 800 44736
rect 1485 44706 1551 44709
rect 0 44704 1551 44706
rect 0 44648 1490 44704
rect 1546 44648 1551 44704
rect 0 44646 1551 44648
rect 0 44616 800 44646
rect 1485 44643 1551 44646
rect 4207 44640 4527 44641
rect 4207 44576 4215 44640
rect 4279 44576 4295 44640
rect 4359 44576 4375 44640
rect 4439 44576 4455 44640
rect 4519 44576 4527 44640
rect 4207 44575 4527 44576
rect 7471 44640 7791 44641
rect 7471 44576 7479 44640
rect 7543 44576 7559 44640
rect 7623 44576 7639 44640
rect 7703 44576 7719 44640
rect 7783 44576 7791 44640
rect 7471 44575 7791 44576
rect 1669 44298 1735 44301
rect 1853 44298 1919 44301
rect 1669 44296 1919 44298
rect 1669 44240 1674 44296
rect 1730 44240 1858 44296
rect 1914 44240 1919 44296
rect 1669 44238 1919 44240
rect 1669 44235 1735 44238
rect 1853 44235 1919 44238
rect 0 44162 800 44192
rect 1577 44162 1643 44165
rect 0 44160 1643 44162
rect 0 44104 1582 44160
rect 1638 44104 1643 44160
rect 0 44102 1643 44104
rect 0 44072 800 44102
rect 1577 44099 1643 44102
rect 2576 44096 2896 44097
rect 2576 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2576 44031 2896 44032
rect 5839 44096 6159 44097
rect 5839 44032 5847 44096
rect 5911 44032 5927 44096
rect 5991 44032 6007 44096
rect 6071 44032 6087 44096
rect 6151 44032 6159 44096
rect 5839 44031 6159 44032
rect 9103 44096 9423 44097
rect 9103 44032 9111 44096
rect 9175 44032 9191 44096
rect 9255 44032 9271 44096
rect 9335 44032 9351 44096
rect 9415 44032 9423 44096
rect 9103 44031 9423 44032
rect 10133 43890 10199 43893
rect 11200 43890 12000 43920
rect 10133 43888 12000 43890
rect 10133 43832 10138 43888
rect 10194 43832 12000 43888
rect 10133 43830 12000 43832
rect 10133 43827 10199 43830
rect 11200 43800 12000 43830
rect 0 43754 800 43784
rect 3969 43754 4035 43757
rect 0 43752 4035 43754
rect 0 43696 3974 43752
rect 4030 43696 4035 43752
rect 0 43694 4035 43696
rect 0 43664 800 43694
rect 3969 43691 4035 43694
rect 4207 43552 4527 43553
rect 4207 43488 4215 43552
rect 4279 43488 4295 43552
rect 4359 43488 4375 43552
rect 4439 43488 4455 43552
rect 4519 43488 4527 43552
rect 4207 43487 4527 43488
rect 7471 43552 7791 43553
rect 7471 43488 7479 43552
rect 7543 43488 7559 43552
rect 7623 43488 7639 43552
rect 7703 43488 7719 43552
rect 7783 43488 7791 43552
rect 7471 43487 7791 43488
rect 0 43346 800 43376
rect 2773 43346 2839 43349
rect 0 43344 2839 43346
rect 0 43288 2778 43344
rect 2834 43288 2839 43344
rect 0 43286 2839 43288
rect 0 43256 800 43286
rect 2773 43283 2839 43286
rect 3141 43210 3207 43213
rect 3734 43210 3740 43212
rect 3141 43208 3740 43210
rect 3141 43152 3146 43208
rect 3202 43152 3740 43208
rect 3141 43150 3740 43152
rect 3141 43147 3207 43150
rect 3734 43148 3740 43150
rect 3804 43148 3810 43212
rect 2576 43008 2896 43009
rect 2576 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2576 42943 2896 42944
rect 5839 43008 6159 43009
rect 5839 42944 5847 43008
rect 5911 42944 5927 43008
rect 5991 42944 6007 43008
rect 6071 42944 6087 43008
rect 6151 42944 6159 43008
rect 5839 42943 6159 42944
rect 9103 43008 9423 43009
rect 9103 42944 9111 43008
rect 9175 42944 9191 43008
rect 9255 42944 9271 43008
rect 9335 42944 9351 43008
rect 9415 42944 9423 43008
rect 9103 42943 9423 42944
rect 0 42802 800 42832
rect 2497 42802 2563 42805
rect 0 42800 2563 42802
rect 0 42744 2502 42800
rect 2558 42744 2563 42800
rect 0 42742 2563 42744
rect 0 42712 800 42742
rect 2497 42739 2563 42742
rect 10041 42802 10107 42805
rect 11200 42802 12000 42832
rect 10041 42800 12000 42802
rect 10041 42744 10046 42800
rect 10102 42744 12000 42800
rect 10041 42742 12000 42744
rect 10041 42739 10107 42742
rect 11200 42712 12000 42742
rect 4207 42464 4527 42465
rect 0 42394 800 42424
rect 4207 42400 4215 42464
rect 4279 42400 4295 42464
rect 4359 42400 4375 42464
rect 4439 42400 4455 42464
rect 4519 42400 4527 42464
rect 4207 42399 4527 42400
rect 7471 42464 7791 42465
rect 7471 42400 7479 42464
rect 7543 42400 7559 42464
rect 7623 42400 7639 42464
rect 7703 42400 7719 42464
rect 7783 42400 7791 42464
rect 7471 42399 7791 42400
rect 2221 42394 2287 42397
rect 0 42392 2287 42394
rect 0 42336 2226 42392
rect 2282 42336 2287 42392
rect 0 42334 2287 42336
rect 0 42304 800 42334
rect 2221 42331 2287 42334
rect 0 41986 800 42016
rect 1485 41986 1551 41989
rect 0 41984 1551 41986
rect 0 41928 1490 41984
rect 1546 41928 1551 41984
rect 0 41926 1551 41928
rect 0 41896 800 41926
rect 1485 41923 1551 41926
rect 2576 41920 2896 41921
rect 2576 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2576 41855 2896 41856
rect 5839 41920 6159 41921
rect 5839 41856 5847 41920
rect 5911 41856 5927 41920
rect 5991 41856 6007 41920
rect 6071 41856 6087 41920
rect 6151 41856 6159 41920
rect 5839 41855 6159 41856
rect 9103 41920 9423 41921
rect 9103 41856 9111 41920
rect 9175 41856 9191 41920
rect 9255 41856 9271 41920
rect 9335 41856 9351 41920
rect 9415 41856 9423 41920
rect 9103 41855 9423 41856
rect 10041 41714 10107 41717
rect 11200 41714 12000 41744
rect 10041 41712 12000 41714
rect 10041 41656 10046 41712
rect 10102 41656 12000 41712
rect 10041 41654 12000 41656
rect 10041 41651 10107 41654
rect 11200 41624 12000 41654
rect 0 41442 800 41472
rect 1393 41442 1459 41445
rect 0 41440 1459 41442
rect 0 41384 1398 41440
rect 1454 41384 1459 41440
rect 0 41382 1459 41384
rect 0 41352 800 41382
rect 1393 41379 1459 41382
rect 4654 41380 4660 41444
rect 4724 41442 4730 41444
rect 5257 41442 5323 41445
rect 4724 41440 5323 41442
rect 4724 41384 5262 41440
rect 5318 41384 5323 41440
rect 4724 41382 5323 41384
rect 4724 41380 4730 41382
rect 5257 41379 5323 41382
rect 4207 41376 4527 41377
rect 4207 41312 4215 41376
rect 4279 41312 4295 41376
rect 4359 41312 4375 41376
rect 4439 41312 4455 41376
rect 4519 41312 4527 41376
rect 4207 41311 4527 41312
rect 7471 41376 7791 41377
rect 7471 41312 7479 41376
rect 7543 41312 7559 41376
rect 7623 41312 7639 41376
rect 7703 41312 7719 41376
rect 7783 41312 7791 41376
rect 7471 41311 7791 41312
rect 0 41034 800 41064
rect 1485 41034 1551 41037
rect 0 41032 1551 41034
rect 0 40976 1490 41032
rect 1546 40976 1551 41032
rect 0 40974 1551 40976
rect 0 40944 800 40974
rect 1485 40971 1551 40974
rect 2576 40832 2896 40833
rect 2576 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2576 40767 2896 40768
rect 5839 40832 6159 40833
rect 5839 40768 5847 40832
rect 5911 40768 5927 40832
rect 5991 40768 6007 40832
rect 6071 40768 6087 40832
rect 6151 40768 6159 40832
rect 5839 40767 6159 40768
rect 9103 40832 9423 40833
rect 9103 40768 9111 40832
rect 9175 40768 9191 40832
rect 9255 40768 9271 40832
rect 9335 40768 9351 40832
rect 9415 40768 9423 40832
rect 9103 40767 9423 40768
rect 0 40626 800 40656
rect 1485 40626 1551 40629
rect 0 40624 1551 40626
rect 0 40568 1490 40624
rect 1546 40568 1551 40624
rect 0 40566 1551 40568
rect 0 40536 800 40566
rect 1485 40563 1551 40566
rect 10041 40626 10107 40629
rect 11200 40626 12000 40656
rect 10041 40624 12000 40626
rect 10041 40568 10046 40624
rect 10102 40568 12000 40624
rect 10041 40566 12000 40568
rect 10041 40563 10107 40566
rect 11200 40536 12000 40566
rect 1669 40354 1735 40357
rect 2078 40354 2084 40356
rect 1669 40352 2084 40354
rect 1669 40296 1674 40352
rect 1730 40296 2084 40352
rect 1669 40294 2084 40296
rect 1669 40291 1735 40294
rect 2078 40292 2084 40294
rect 2148 40292 2154 40356
rect 4207 40288 4527 40289
rect 0 40218 800 40248
rect 4207 40224 4215 40288
rect 4279 40224 4295 40288
rect 4359 40224 4375 40288
rect 4439 40224 4455 40288
rect 4519 40224 4527 40288
rect 4207 40223 4527 40224
rect 7471 40288 7791 40289
rect 7471 40224 7479 40288
rect 7543 40224 7559 40288
rect 7623 40224 7639 40288
rect 7703 40224 7719 40288
rect 7783 40224 7791 40288
rect 7471 40223 7791 40224
rect 1485 40218 1551 40221
rect 0 40216 1551 40218
rect 0 40160 1490 40216
rect 1546 40160 1551 40216
rect 0 40158 1551 40160
rect 0 40128 800 40158
rect 1485 40155 1551 40158
rect 1853 40082 1919 40085
rect 2262 40082 2268 40084
rect 1853 40080 2268 40082
rect 1853 40024 1858 40080
rect 1914 40024 2268 40080
rect 1853 40022 2268 40024
rect 1853 40019 1919 40022
rect 2262 40020 2268 40022
rect 2332 40020 2338 40084
rect 2576 39744 2896 39745
rect 0 39674 800 39704
rect 2576 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2576 39679 2896 39680
rect 5839 39744 6159 39745
rect 5839 39680 5847 39744
rect 5911 39680 5927 39744
rect 5991 39680 6007 39744
rect 6071 39680 6087 39744
rect 6151 39680 6159 39744
rect 5839 39679 6159 39680
rect 9103 39744 9423 39745
rect 9103 39680 9111 39744
rect 9175 39680 9191 39744
rect 9255 39680 9271 39744
rect 9335 39680 9351 39744
rect 9415 39680 9423 39744
rect 9103 39679 9423 39680
rect 1485 39674 1551 39677
rect 0 39672 1551 39674
rect 0 39616 1490 39672
rect 1546 39616 1551 39672
rect 0 39614 1551 39616
rect 0 39584 800 39614
rect 1485 39611 1551 39614
rect 10041 39402 10107 39405
rect 11200 39402 12000 39432
rect 10041 39400 12000 39402
rect 10041 39344 10046 39400
rect 10102 39344 12000 39400
rect 10041 39342 12000 39344
rect 10041 39339 10107 39342
rect 11200 39312 12000 39342
rect 0 39266 800 39296
rect 1485 39266 1551 39269
rect 0 39264 1551 39266
rect 0 39208 1490 39264
rect 1546 39208 1551 39264
rect 0 39206 1551 39208
rect 0 39176 800 39206
rect 1485 39203 1551 39206
rect 4207 39200 4527 39201
rect 4207 39136 4215 39200
rect 4279 39136 4295 39200
rect 4359 39136 4375 39200
rect 4439 39136 4455 39200
rect 4519 39136 4527 39200
rect 4207 39135 4527 39136
rect 7471 39200 7791 39201
rect 7471 39136 7479 39200
rect 7543 39136 7559 39200
rect 7623 39136 7639 39200
rect 7703 39136 7719 39200
rect 7783 39136 7791 39200
rect 7471 39135 7791 39136
rect 0 38858 800 38888
rect 1485 38858 1551 38861
rect 0 38856 1551 38858
rect 0 38800 1490 38856
rect 1546 38800 1551 38856
rect 0 38798 1551 38800
rect 0 38768 800 38798
rect 1485 38795 1551 38798
rect 2576 38656 2896 38657
rect 2576 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2576 38591 2896 38592
rect 5839 38656 6159 38657
rect 5839 38592 5847 38656
rect 5911 38592 5927 38656
rect 5991 38592 6007 38656
rect 6071 38592 6087 38656
rect 6151 38592 6159 38656
rect 5839 38591 6159 38592
rect 9103 38656 9423 38657
rect 9103 38592 9111 38656
rect 9175 38592 9191 38656
rect 9255 38592 9271 38656
rect 9335 38592 9351 38656
rect 9415 38592 9423 38656
rect 9103 38591 9423 38592
rect 0 38314 800 38344
rect 1393 38314 1459 38317
rect 0 38312 1459 38314
rect 0 38256 1398 38312
rect 1454 38256 1459 38312
rect 0 38254 1459 38256
rect 0 38224 800 38254
rect 1393 38251 1459 38254
rect 10041 38314 10107 38317
rect 11200 38314 12000 38344
rect 10041 38312 12000 38314
rect 10041 38256 10046 38312
rect 10102 38256 12000 38312
rect 10041 38254 12000 38256
rect 10041 38251 10107 38254
rect 11200 38224 12000 38254
rect 4207 38112 4527 38113
rect 4207 38048 4215 38112
rect 4279 38048 4295 38112
rect 4359 38048 4375 38112
rect 4439 38048 4455 38112
rect 4519 38048 4527 38112
rect 4207 38047 4527 38048
rect 7471 38112 7791 38113
rect 7471 38048 7479 38112
rect 7543 38048 7559 38112
rect 7623 38048 7639 38112
rect 7703 38048 7719 38112
rect 7783 38048 7791 38112
rect 7471 38047 7791 38048
rect 0 37906 800 37936
rect 1485 37906 1551 37909
rect 0 37904 1551 37906
rect 0 37848 1490 37904
rect 1546 37848 1551 37904
rect 0 37846 1551 37848
rect 0 37816 800 37846
rect 1485 37843 1551 37846
rect 2576 37568 2896 37569
rect 0 37498 800 37528
rect 2576 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2576 37503 2896 37504
rect 5839 37568 6159 37569
rect 5839 37504 5847 37568
rect 5911 37504 5927 37568
rect 5991 37504 6007 37568
rect 6071 37504 6087 37568
rect 6151 37504 6159 37568
rect 5839 37503 6159 37504
rect 9103 37568 9423 37569
rect 9103 37504 9111 37568
rect 9175 37504 9191 37568
rect 9255 37504 9271 37568
rect 9335 37504 9351 37568
rect 9415 37504 9423 37568
rect 9103 37503 9423 37504
rect 0 37438 1778 37498
rect 0 37408 800 37438
rect 1718 37362 1778 37438
rect 3233 37362 3299 37365
rect 1718 37360 3299 37362
rect 1718 37304 3238 37360
rect 3294 37304 3299 37360
rect 1718 37302 3299 37304
rect 3233 37299 3299 37302
rect 10041 37226 10107 37229
rect 11200 37226 12000 37256
rect 10041 37224 12000 37226
rect 10041 37168 10046 37224
rect 10102 37168 12000 37224
rect 10041 37166 12000 37168
rect 10041 37163 10107 37166
rect 11200 37136 12000 37166
rect 4207 37024 4527 37025
rect 0 36954 800 36984
rect 4207 36960 4215 37024
rect 4279 36960 4295 37024
rect 4359 36960 4375 37024
rect 4439 36960 4455 37024
rect 4519 36960 4527 37024
rect 4207 36959 4527 36960
rect 7471 37024 7791 37025
rect 7471 36960 7479 37024
rect 7543 36960 7559 37024
rect 7623 36960 7639 37024
rect 7703 36960 7719 37024
rect 7783 36960 7791 37024
rect 7471 36959 7791 36960
rect 2313 36954 2379 36957
rect 0 36952 2379 36954
rect 0 36896 2318 36952
rect 2374 36896 2379 36952
rect 0 36894 2379 36896
rect 0 36864 800 36894
rect 2313 36891 2379 36894
rect 2078 36756 2084 36820
rect 2148 36818 2154 36820
rect 2313 36818 2379 36821
rect 2148 36816 2379 36818
rect 2148 36760 2318 36816
rect 2374 36760 2379 36816
rect 2148 36758 2379 36760
rect 2148 36756 2154 36758
rect 2313 36755 2379 36758
rect 0 36546 800 36576
rect 1577 36546 1643 36549
rect 0 36544 1643 36546
rect 0 36488 1582 36544
rect 1638 36488 1643 36544
rect 0 36486 1643 36488
rect 0 36456 800 36486
rect 1577 36483 1643 36486
rect 2576 36480 2896 36481
rect 2576 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2576 36415 2896 36416
rect 5839 36480 6159 36481
rect 5839 36416 5847 36480
rect 5911 36416 5927 36480
rect 5991 36416 6007 36480
rect 6071 36416 6087 36480
rect 6151 36416 6159 36480
rect 5839 36415 6159 36416
rect 9103 36480 9423 36481
rect 9103 36416 9111 36480
rect 9175 36416 9191 36480
rect 9255 36416 9271 36480
rect 9335 36416 9351 36480
rect 9415 36416 9423 36480
rect 9103 36415 9423 36416
rect 0 36138 800 36168
rect 1485 36138 1551 36141
rect 0 36136 1551 36138
rect 0 36080 1490 36136
rect 1546 36080 1551 36136
rect 0 36078 1551 36080
rect 0 36048 800 36078
rect 1485 36075 1551 36078
rect 10041 36138 10107 36141
rect 11200 36138 12000 36168
rect 10041 36136 12000 36138
rect 10041 36080 10046 36136
rect 10102 36080 12000 36136
rect 10041 36078 12000 36080
rect 10041 36075 10107 36078
rect 11200 36048 12000 36078
rect 4207 35936 4527 35937
rect 4207 35872 4215 35936
rect 4279 35872 4295 35936
rect 4359 35872 4375 35936
rect 4439 35872 4455 35936
rect 4519 35872 4527 35936
rect 4207 35871 4527 35872
rect 7471 35936 7791 35937
rect 7471 35872 7479 35936
rect 7543 35872 7559 35936
rect 7623 35872 7639 35936
rect 7703 35872 7719 35936
rect 7783 35872 7791 35936
rect 7471 35871 7791 35872
rect 2129 35866 2195 35869
rect 2589 35866 2655 35869
rect 2129 35864 2655 35866
rect 2129 35808 2134 35864
rect 2190 35808 2594 35864
rect 2650 35808 2655 35864
rect 2129 35806 2655 35808
rect 2129 35803 2195 35806
rect 2589 35803 2655 35806
rect 0 35594 800 35624
rect 2313 35594 2379 35597
rect 0 35592 2379 35594
rect 0 35536 2318 35592
rect 2374 35536 2379 35592
rect 0 35534 2379 35536
rect 0 35504 800 35534
rect 2313 35531 2379 35534
rect 2576 35392 2896 35393
rect 2576 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2576 35327 2896 35328
rect 5839 35392 6159 35393
rect 5839 35328 5847 35392
rect 5911 35328 5927 35392
rect 5991 35328 6007 35392
rect 6071 35328 6087 35392
rect 6151 35328 6159 35392
rect 5839 35327 6159 35328
rect 9103 35392 9423 35393
rect 9103 35328 9111 35392
rect 9175 35328 9191 35392
rect 9255 35328 9271 35392
rect 9335 35328 9351 35392
rect 9415 35328 9423 35392
rect 9103 35327 9423 35328
rect 0 35186 800 35216
rect 1577 35186 1643 35189
rect 0 35184 1643 35186
rect 0 35128 1582 35184
rect 1638 35128 1643 35184
rect 0 35126 1643 35128
rect 0 35096 800 35126
rect 1577 35123 1643 35126
rect 10041 35050 10107 35053
rect 11200 35050 12000 35080
rect 10041 35048 12000 35050
rect 10041 34992 10046 35048
rect 10102 34992 12000 35048
rect 10041 34990 12000 34992
rect 10041 34987 10107 34990
rect 11200 34960 12000 34990
rect 4207 34848 4527 34849
rect 0 34778 800 34808
rect 4207 34784 4215 34848
rect 4279 34784 4295 34848
rect 4359 34784 4375 34848
rect 4439 34784 4455 34848
rect 4519 34784 4527 34848
rect 4207 34783 4527 34784
rect 7471 34848 7791 34849
rect 7471 34784 7479 34848
rect 7543 34784 7559 34848
rect 7623 34784 7639 34848
rect 7703 34784 7719 34848
rect 7783 34784 7791 34848
rect 7471 34783 7791 34784
rect 1485 34778 1551 34781
rect 0 34776 1551 34778
rect 0 34720 1490 34776
rect 1546 34720 1551 34776
rect 0 34718 1551 34720
rect 0 34688 800 34718
rect 1485 34715 1551 34718
rect 0 34370 800 34400
rect 1577 34370 1643 34373
rect 0 34368 1643 34370
rect 0 34312 1582 34368
rect 1638 34312 1643 34368
rect 0 34310 1643 34312
rect 0 34280 800 34310
rect 1577 34307 1643 34310
rect 2576 34304 2896 34305
rect 2576 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2576 34239 2896 34240
rect 5839 34304 6159 34305
rect 5839 34240 5847 34304
rect 5911 34240 5927 34304
rect 5991 34240 6007 34304
rect 6071 34240 6087 34304
rect 6151 34240 6159 34304
rect 5839 34239 6159 34240
rect 9103 34304 9423 34305
rect 9103 34240 9111 34304
rect 9175 34240 9191 34304
rect 9255 34240 9271 34304
rect 9335 34240 9351 34304
rect 9415 34240 9423 34304
rect 9103 34239 9423 34240
rect 10041 33962 10107 33965
rect 11200 33962 12000 33992
rect 10041 33960 12000 33962
rect 10041 33904 10046 33960
rect 10102 33904 12000 33960
rect 10041 33902 12000 33904
rect 10041 33899 10107 33902
rect 11200 33872 12000 33902
rect 0 33826 800 33856
rect 1485 33826 1551 33829
rect 0 33824 1551 33826
rect 0 33768 1490 33824
rect 1546 33768 1551 33824
rect 0 33766 1551 33768
rect 0 33736 800 33766
rect 1485 33763 1551 33766
rect 4207 33760 4527 33761
rect 4207 33696 4215 33760
rect 4279 33696 4295 33760
rect 4359 33696 4375 33760
rect 4439 33696 4455 33760
rect 4519 33696 4527 33760
rect 4207 33695 4527 33696
rect 7471 33760 7791 33761
rect 7471 33696 7479 33760
rect 7543 33696 7559 33760
rect 7623 33696 7639 33760
rect 7703 33696 7719 33760
rect 7783 33696 7791 33760
rect 7471 33695 7791 33696
rect 0 33418 800 33448
rect 1577 33418 1643 33421
rect 0 33416 1643 33418
rect 0 33360 1582 33416
rect 1638 33360 1643 33416
rect 0 33358 1643 33360
rect 0 33328 800 33358
rect 1577 33355 1643 33358
rect 2576 33216 2896 33217
rect 2576 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2576 33151 2896 33152
rect 5839 33216 6159 33217
rect 5839 33152 5847 33216
rect 5911 33152 5927 33216
rect 5991 33152 6007 33216
rect 6071 33152 6087 33216
rect 6151 33152 6159 33216
rect 5839 33151 6159 33152
rect 9103 33216 9423 33217
rect 9103 33152 9111 33216
rect 9175 33152 9191 33216
rect 9255 33152 9271 33216
rect 9335 33152 9351 33216
rect 9415 33152 9423 33216
rect 9103 33151 9423 33152
rect 0 33010 800 33040
rect 1577 33010 1643 33013
rect 0 33008 1643 33010
rect 0 32952 1582 33008
rect 1638 32952 1643 33008
rect 0 32950 1643 32952
rect 0 32920 800 32950
rect 1577 32947 1643 32950
rect 10041 32738 10107 32741
rect 11200 32738 12000 32768
rect 10041 32736 12000 32738
rect 10041 32680 10046 32736
rect 10102 32680 12000 32736
rect 10041 32678 12000 32680
rect 10041 32675 10107 32678
rect 4207 32672 4527 32673
rect 4207 32608 4215 32672
rect 4279 32608 4295 32672
rect 4359 32608 4375 32672
rect 4439 32608 4455 32672
rect 4519 32608 4527 32672
rect 4207 32607 4527 32608
rect 7471 32672 7791 32673
rect 7471 32608 7479 32672
rect 7543 32608 7559 32672
rect 7623 32608 7639 32672
rect 7703 32608 7719 32672
rect 7783 32608 7791 32672
rect 11200 32648 12000 32678
rect 7471 32607 7791 32608
rect 0 32466 800 32496
rect 3049 32466 3115 32469
rect 0 32464 3115 32466
rect 0 32408 3054 32464
rect 3110 32408 3115 32464
rect 0 32406 3115 32408
rect 0 32376 800 32406
rect 3049 32403 3115 32406
rect 3233 32330 3299 32333
rect 1718 32328 3299 32330
rect 1718 32272 3238 32328
rect 3294 32272 3299 32328
rect 1718 32270 3299 32272
rect 0 32058 800 32088
rect 1718 32058 1778 32270
rect 3233 32267 3299 32270
rect 2576 32128 2896 32129
rect 2576 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2576 32063 2896 32064
rect 5839 32128 6159 32129
rect 5839 32064 5847 32128
rect 5911 32064 5927 32128
rect 5991 32064 6007 32128
rect 6071 32064 6087 32128
rect 6151 32064 6159 32128
rect 5839 32063 6159 32064
rect 9103 32128 9423 32129
rect 9103 32064 9111 32128
rect 9175 32064 9191 32128
rect 9255 32064 9271 32128
rect 9335 32064 9351 32128
rect 9415 32064 9423 32128
rect 9103 32063 9423 32064
rect 0 31998 1778 32058
rect 0 31968 800 31998
rect 0 31650 800 31680
rect 2773 31650 2839 31653
rect 0 31648 2839 31650
rect 0 31592 2778 31648
rect 2834 31592 2839 31648
rect 0 31590 2839 31592
rect 0 31560 800 31590
rect 2773 31587 2839 31590
rect 10041 31650 10107 31653
rect 11200 31650 12000 31680
rect 10041 31648 12000 31650
rect 10041 31592 10046 31648
rect 10102 31592 12000 31648
rect 10041 31590 12000 31592
rect 10041 31587 10107 31590
rect 4207 31584 4527 31585
rect 4207 31520 4215 31584
rect 4279 31520 4295 31584
rect 4359 31520 4375 31584
rect 4439 31520 4455 31584
rect 4519 31520 4527 31584
rect 4207 31519 4527 31520
rect 7471 31584 7791 31585
rect 7471 31520 7479 31584
rect 7543 31520 7559 31584
rect 7623 31520 7639 31584
rect 7703 31520 7719 31584
rect 7783 31520 7791 31584
rect 11200 31560 12000 31590
rect 7471 31519 7791 31520
rect 0 31106 800 31136
rect 1393 31106 1459 31109
rect 0 31104 1459 31106
rect 0 31048 1398 31104
rect 1454 31048 1459 31104
rect 0 31046 1459 31048
rect 0 31016 800 31046
rect 1393 31043 1459 31046
rect 2576 31040 2896 31041
rect 2576 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2576 30975 2896 30976
rect 5839 31040 6159 31041
rect 5839 30976 5847 31040
rect 5911 30976 5927 31040
rect 5991 30976 6007 31040
rect 6071 30976 6087 31040
rect 6151 30976 6159 31040
rect 5839 30975 6159 30976
rect 9103 31040 9423 31041
rect 9103 30976 9111 31040
rect 9175 30976 9191 31040
rect 9255 30976 9271 31040
rect 9335 30976 9351 31040
rect 9415 30976 9423 31040
rect 9103 30975 9423 30976
rect 0 30698 800 30728
rect 3969 30698 4035 30701
rect 0 30696 4035 30698
rect 0 30640 3974 30696
rect 4030 30640 4035 30696
rect 0 30638 4035 30640
rect 0 30608 800 30638
rect 3969 30635 4035 30638
rect 10041 30562 10107 30565
rect 11200 30562 12000 30592
rect 10041 30560 12000 30562
rect 10041 30504 10046 30560
rect 10102 30504 12000 30560
rect 10041 30502 12000 30504
rect 10041 30499 10107 30502
rect 4207 30496 4527 30497
rect 4207 30432 4215 30496
rect 4279 30432 4295 30496
rect 4359 30432 4375 30496
rect 4439 30432 4455 30496
rect 4519 30432 4527 30496
rect 4207 30431 4527 30432
rect 7471 30496 7791 30497
rect 7471 30432 7479 30496
rect 7543 30432 7559 30496
rect 7623 30432 7639 30496
rect 7703 30432 7719 30496
rect 7783 30432 7791 30496
rect 11200 30472 12000 30502
rect 7471 30431 7791 30432
rect 0 30290 800 30320
rect 3141 30290 3207 30293
rect 0 30288 3207 30290
rect 0 30232 3146 30288
rect 3202 30232 3207 30288
rect 0 30230 3207 30232
rect 0 30200 800 30230
rect 3141 30227 3207 30230
rect 2773 30154 2839 30157
rect 1350 30152 2839 30154
rect 1350 30096 2778 30152
rect 2834 30096 2839 30152
rect 1350 30094 2839 30096
rect 0 29882 800 29912
rect 1350 29882 1410 30094
rect 2773 30091 2839 30094
rect 2576 29952 2896 29953
rect 2576 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2576 29887 2896 29888
rect 5839 29952 6159 29953
rect 5839 29888 5847 29952
rect 5911 29888 5927 29952
rect 5991 29888 6007 29952
rect 6071 29888 6087 29952
rect 6151 29888 6159 29952
rect 5839 29887 6159 29888
rect 9103 29952 9423 29953
rect 9103 29888 9111 29952
rect 9175 29888 9191 29952
rect 9255 29888 9271 29952
rect 9335 29888 9351 29952
rect 9415 29888 9423 29952
rect 9103 29887 9423 29888
rect 0 29822 1410 29882
rect 0 29792 800 29822
rect 10041 29474 10107 29477
rect 11200 29474 12000 29504
rect 10041 29472 12000 29474
rect 10041 29416 10046 29472
rect 10102 29416 12000 29472
rect 10041 29414 12000 29416
rect 10041 29411 10107 29414
rect 4207 29408 4527 29409
rect 0 29338 800 29368
rect 4207 29344 4215 29408
rect 4279 29344 4295 29408
rect 4359 29344 4375 29408
rect 4439 29344 4455 29408
rect 4519 29344 4527 29408
rect 4207 29343 4527 29344
rect 7471 29408 7791 29409
rect 7471 29344 7479 29408
rect 7543 29344 7559 29408
rect 7623 29344 7639 29408
rect 7703 29344 7719 29408
rect 7783 29344 7791 29408
rect 11200 29384 12000 29414
rect 7471 29343 7791 29344
rect 3233 29338 3299 29341
rect 0 29336 3299 29338
rect 0 29280 3238 29336
rect 3294 29280 3299 29336
rect 0 29278 3299 29280
rect 0 29248 800 29278
rect 3233 29275 3299 29278
rect 0 28930 800 28960
rect 2313 28930 2379 28933
rect 0 28928 2379 28930
rect 0 28872 2318 28928
rect 2374 28872 2379 28928
rect 0 28870 2379 28872
rect 0 28840 800 28870
rect 2313 28867 2379 28870
rect 2576 28864 2896 28865
rect 2576 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2576 28799 2896 28800
rect 5839 28864 6159 28865
rect 5839 28800 5847 28864
rect 5911 28800 5927 28864
rect 5991 28800 6007 28864
rect 6071 28800 6087 28864
rect 6151 28800 6159 28864
rect 5839 28799 6159 28800
rect 9103 28864 9423 28865
rect 9103 28800 9111 28864
rect 9175 28800 9191 28864
rect 9255 28800 9271 28864
rect 9335 28800 9351 28864
rect 9415 28800 9423 28864
rect 9103 28799 9423 28800
rect 0 28522 800 28552
rect 3509 28522 3575 28525
rect 0 28520 3575 28522
rect 0 28464 3514 28520
rect 3570 28464 3575 28520
rect 0 28462 3575 28464
rect 0 28432 800 28462
rect 3509 28459 3575 28462
rect 10041 28386 10107 28389
rect 11200 28386 12000 28416
rect 10041 28384 12000 28386
rect 10041 28328 10046 28384
rect 10102 28328 12000 28384
rect 10041 28326 12000 28328
rect 10041 28323 10107 28326
rect 4207 28320 4527 28321
rect 4207 28256 4215 28320
rect 4279 28256 4295 28320
rect 4359 28256 4375 28320
rect 4439 28256 4455 28320
rect 4519 28256 4527 28320
rect 4207 28255 4527 28256
rect 7471 28320 7791 28321
rect 7471 28256 7479 28320
rect 7543 28256 7559 28320
rect 7623 28256 7639 28320
rect 7703 28256 7719 28320
rect 7783 28256 7791 28320
rect 11200 28296 12000 28326
rect 7471 28255 7791 28256
rect 0 27978 800 28008
rect 3049 27978 3115 27981
rect 0 27976 3115 27978
rect 0 27920 3054 27976
rect 3110 27920 3115 27976
rect 0 27918 3115 27920
rect 0 27888 800 27918
rect 3049 27915 3115 27918
rect 2576 27776 2896 27777
rect 2576 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2576 27711 2896 27712
rect 5839 27776 6159 27777
rect 5839 27712 5847 27776
rect 5911 27712 5927 27776
rect 5991 27712 6007 27776
rect 6071 27712 6087 27776
rect 6151 27712 6159 27776
rect 5839 27711 6159 27712
rect 9103 27776 9423 27777
rect 9103 27712 9111 27776
rect 9175 27712 9191 27776
rect 9255 27712 9271 27776
rect 9335 27712 9351 27776
rect 9415 27712 9423 27776
rect 9103 27711 9423 27712
rect 0 27570 800 27600
rect 3141 27570 3207 27573
rect 0 27568 3207 27570
rect 0 27512 3146 27568
rect 3202 27512 3207 27568
rect 0 27510 3207 27512
rect 0 27480 800 27510
rect 3141 27507 3207 27510
rect 10041 27298 10107 27301
rect 11200 27298 12000 27328
rect 10041 27296 12000 27298
rect 10041 27240 10046 27296
rect 10102 27240 12000 27296
rect 10041 27238 12000 27240
rect 10041 27235 10107 27238
rect 4207 27232 4527 27233
rect 0 27162 800 27192
rect 4207 27168 4215 27232
rect 4279 27168 4295 27232
rect 4359 27168 4375 27232
rect 4439 27168 4455 27232
rect 4519 27168 4527 27232
rect 4207 27167 4527 27168
rect 7471 27232 7791 27233
rect 7471 27168 7479 27232
rect 7543 27168 7559 27232
rect 7623 27168 7639 27232
rect 7703 27168 7719 27232
rect 7783 27168 7791 27232
rect 11200 27208 12000 27238
rect 7471 27167 7791 27168
rect 2221 27162 2287 27165
rect 0 27160 2287 27162
rect 0 27104 2226 27160
rect 2282 27104 2287 27160
rect 0 27102 2287 27104
rect 0 27072 800 27102
rect 2221 27099 2287 27102
rect 2865 26890 2931 26893
rect 1488 26888 2931 26890
rect 1488 26832 2870 26888
rect 2926 26832 2931 26888
rect 1488 26830 2931 26832
rect 0 26618 800 26648
rect 1488 26618 1548 26830
rect 2865 26827 2931 26830
rect 2576 26688 2896 26689
rect 2576 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2576 26623 2896 26624
rect 5839 26688 6159 26689
rect 5839 26624 5847 26688
rect 5911 26624 5927 26688
rect 5991 26624 6007 26688
rect 6071 26624 6087 26688
rect 6151 26624 6159 26688
rect 5839 26623 6159 26624
rect 9103 26688 9423 26689
rect 9103 26624 9111 26688
rect 9175 26624 9191 26688
rect 9255 26624 9271 26688
rect 9335 26624 9351 26688
rect 9415 26624 9423 26688
rect 9103 26623 9423 26624
rect 0 26558 1548 26618
rect 0 26528 800 26558
rect 0 26210 800 26240
rect 2037 26210 2103 26213
rect 0 26208 2103 26210
rect 0 26152 2042 26208
rect 2098 26152 2103 26208
rect 0 26150 2103 26152
rect 0 26120 800 26150
rect 2037 26147 2103 26150
rect 4207 26144 4527 26145
rect 4207 26080 4215 26144
rect 4279 26080 4295 26144
rect 4359 26080 4375 26144
rect 4439 26080 4455 26144
rect 4519 26080 4527 26144
rect 4207 26079 4527 26080
rect 7471 26144 7791 26145
rect 7471 26080 7479 26144
rect 7543 26080 7559 26144
rect 7623 26080 7639 26144
rect 7703 26080 7719 26144
rect 7783 26080 7791 26144
rect 7471 26079 7791 26080
rect 10041 26074 10107 26077
rect 11200 26074 12000 26104
rect 10041 26072 12000 26074
rect 10041 26016 10046 26072
rect 10102 26016 12000 26072
rect 10041 26014 12000 26016
rect 10041 26011 10107 26014
rect 11200 25984 12000 26014
rect 0 25802 800 25832
rect 2221 25802 2287 25805
rect 0 25800 2287 25802
rect 0 25744 2226 25800
rect 2282 25744 2287 25800
rect 0 25742 2287 25744
rect 0 25712 800 25742
rect 2221 25739 2287 25742
rect 2576 25600 2896 25601
rect 2576 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2576 25535 2896 25536
rect 5839 25600 6159 25601
rect 5839 25536 5847 25600
rect 5911 25536 5927 25600
rect 5991 25536 6007 25600
rect 6071 25536 6087 25600
rect 6151 25536 6159 25600
rect 5839 25535 6159 25536
rect 9103 25600 9423 25601
rect 9103 25536 9111 25600
rect 9175 25536 9191 25600
rect 9255 25536 9271 25600
rect 9335 25536 9351 25600
rect 9415 25536 9423 25600
rect 9103 25535 9423 25536
rect 0 25258 800 25288
rect 2865 25258 2931 25261
rect 0 25256 2931 25258
rect 0 25200 2870 25256
rect 2926 25200 2931 25256
rect 0 25198 2931 25200
rect 0 25168 800 25198
rect 2865 25195 2931 25198
rect 4207 25056 4527 25057
rect 4207 24992 4215 25056
rect 4279 24992 4295 25056
rect 4359 24992 4375 25056
rect 4439 24992 4455 25056
rect 4519 24992 4527 25056
rect 4207 24991 4527 24992
rect 7471 25056 7791 25057
rect 7471 24992 7479 25056
rect 7543 24992 7559 25056
rect 7623 24992 7639 25056
rect 7703 24992 7719 25056
rect 7783 24992 7791 25056
rect 7471 24991 7791 24992
rect 10041 24986 10107 24989
rect 11200 24986 12000 25016
rect 10041 24984 12000 24986
rect 10041 24928 10046 24984
rect 10102 24928 12000 24984
rect 10041 24926 12000 24928
rect 10041 24923 10107 24926
rect 11200 24896 12000 24926
rect 0 24850 800 24880
rect 2221 24850 2287 24853
rect 0 24848 2287 24850
rect 0 24792 2226 24848
rect 2282 24792 2287 24848
rect 0 24790 2287 24792
rect 0 24760 800 24790
rect 2221 24787 2287 24790
rect 1393 24712 1459 24717
rect 1393 24656 1398 24712
rect 1454 24656 1459 24712
rect 1393 24651 1459 24656
rect 0 24442 800 24472
rect 1396 24442 1456 24651
rect 2576 24512 2896 24513
rect 2576 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2576 24447 2896 24448
rect 5839 24512 6159 24513
rect 5839 24448 5847 24512
rect 5911 24448 5927 24512
rect 5991 24448 6007 24512
rect 6071 24448 6087 24512
rect 6151 24448 6159 24512
rect 5839 24447 6159 24448
rect 9103 24512 9423 24513
rect 9103 24448 9111 24512
rect 9175 24448 9191 24512
rect 9255 24448 9271 24512
rect 9335 24448 9351 24512
rect 9415 24448 9423 24512
rect 9103 24447 9423 24448
rect 0 24382 1456 24442
rect 0 24352 800 24382
rect 0 24034 800 24064
rect 2865 24034 2931 24037
rect 0 24032 2931 24034
rect 0 23976 2870 24032
rect 2926 23976 2931 24032
rect 0 23974 2931 23976
rect 0 23944 800 23974
rect 2865 23971 2931 23974
rect 4207 23968 4527 23969
rect 4207 23904 4215 23968
rect 4279 23904 4295 23968
rect 4359 23904 4375 23968
rect 4439 23904 4455 23968
rect 4519 23904 4527 23968
rect 4207 23903 4527 23904
rect 7471 23968 7791 23969
rect 7471 23904 7479 23968
rect 7543 23904 7559 23968
rect 7623 23904 7639 23968
rect 7703 23904 7719 23968
rect 7783 23904 7791 23968
rect 7471 23903 7791 23904
rect 10041 23898 10107 23901
rect 11200 23898 12000 23928
rect 10041 23896 12000 23898
rect 10041 23840 10046 23896
rect 10102 23840 12000 23896
rect 10041 23838 12000 23840
rect 10041 23835 10107 23838
rect 11200 23808 12000 23838
rect 1158 23564 1164 23628
rect 1228 23626 1234 23628
rect 2037 23626 2103 23629
rect 1228 23624 2103 23626
rect 1228 23568 2042 23624
rect 2098 23568 2103 23624
rect 1228 23566 2103 23568
rect 1228 23564 1234 23566
rect 2037 23563 2103 23566
rect 0 23490 800 23520
rect 1485 23490 1551 23493
rect 0 23488 1551 23490
rect 0 23432 1490 23488
rect 1546 23432 1551 23488
rect 0 23430 1551 23432
rect 0 23400 800 23430
rect 1485 23427 1551 23430
rect 2576 23424 2896 23425
rect 2576 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2576 23359 2896 23360
rect 5839 23424 6159 23425
rect 5839 23360 5847 23424
rect 5911 23360 5927 23424
rect 5991 23360 6007 23424
rect 6071 23360 6087 23424
rect 6151 23360 6159 23424
rect 5839 23359 6159 23360
rect 9103 23424 9423 23425
rect 9103 23360 9111 23424
rect 9175 23360 9191 23424
rect 9255 23360 9271 23424
rect 9335 23360 9351 23424
rect 9415 23360 9423 23424
rect 9103 23359 9423 23360
rect 0 23082 800 23112
rect 1485 23082 1551 23085
rect 0 23080 1551 23082
rect 0 23024 1490 23080
rect 1546 23024 1551 23080
rect 0 23022 1551 23024
rect 0 22992 800 23022
rect 1485 23019 1551 23022
rect 4207 22880 4527 22881
rect 4207 22816 4215 22880
rect 4279 22816 4295 22880
rect 4359 22816 4375 22880
rect 4439 22816 4455 22880
rect 4519 22816 4527 22880
rect 4207 22815 4527 22816
rect 7471 22880 7791 22881
rect 7471 22816 7479 22880
rect 7543 22816 7559 22880
rect 7623 22816 7639 22880
rect 7703 22816 7719 22880
rect 7783 22816 7791 22880
rect 7471 22815 7791 22816
rect 10041 22810 10107 22813
rect 11200 22810 12000 22840
rect 10041 22808 12000 22810
rect 10041 22752 10046 22808
rect 10102 22752 12000 22808
rect 10041 22750 12000 22752
rect 10041 22747 10107 22750
rect 11200 22720 12000 22750
rect 0 22674 800 22704
rect 3785 22674 3851 22677
rect 0 22672 3851 22674
rect 0 22616 3790 22672
rect 3846 22616 3851 22672
rect 0 22614 3851 22616
rect 0 22584 800 22614
rect 3785 22611 3851 22614
rect 2576 22336 2896 22337
rect 2576 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2576 22271 2896 22272
rect 5839 22336 6159 22337
rect 5839 22272 5847 22336
rect 5911 22272 5927 22336
rect 5991 22272 6007 22336
rect 6071 22272 6087 22336
rect 6151 22272 6159 22336
rect 5839 22271 6159 22272
rect 9103 22336 9423 22337
rect 9103 22272 9111 22336
rect 9175 22272 9191 22336
rect 9255 22272 9271 22336
rect 9335 22272 9351 22336
rect 9415 22272 9423 22336
rect 9103 22271 9423 22272
rect 0 22130 800 22160
rect 3325 22130 3391 22133
rect 0 22128 3391 22130
rect 0 22072 3330 22128
rect 3386 22072 3391 22128
rect 0 22070 3391 22072
rect 0 22040 800 22070
rect 3325 22067 3391 22070
rect 4207 21792 4527 21793
rect 0 21722 800 21752
rect 4207 21728 4215 21792
rect 4279 21728 4295 21792
rect 4359 21728 4375 21792
rect 4439 21728 4455 21792
rect 4519 21728 4527 21792
rect 4207 21727 4527 21728
rect 7471 21792 7791 21793
rect 7471 21728 7479 21792
rect 7543 21728 7559 21792
rect 7623 21728 7639 21792
rect 7703 21728 7719 21792
rect 7783 21728 7791 21792
rect 7471 21727 7791 21728
rect 2037 21722 2103 21725
rect 0 21720 2103 21722
rect 0 21664 2042 21720
rect 2098 21664 2103 21720
rect 0 21662 2103 21664
rect 0 21632 800 21662
rect 2037 21659 2103 21662
rect 10041 21722 10107 21725
rect 11200 21722 12000 21752
rect 10041 21720 12000 21722
rect 10041 21664 10046 21720
rect 10102 21664 12000 21720
rect 10041 21662 12000 21664
rect 10041 21659 10107 21662
rect 11200 21632 12000 21662
rect 2865 21450 2931 21453
rect 1396 21448 2931 21450
rect 1396 21392 2870 21448
rect 2926 21392 2931 21448
rect 1396 21390 2931 21392
rect 0 21314 800 21344
rect 1396 21314 1456 21390
rect 2865 21387 2931 21390
rect 0 21254 1456 21314
rect 0 21224 800 21254
rect 2576 21248 2896 21249
rect 2576 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2576 21183 2896 21184
rect 5839 21248 6159 21249
rect 5839 21184 5847 21248
rect 5911 21184 5927 21248
rect 5991 21184 6007 21248
rect 6071 21184 6087 21248
rect 6151 21184 6159 21248
rect 5839 21183 6159 21184
rect 9103 21248 9423 21249
rect 9103 21184 9111 21248
rect 9175 21184 9191 21248
rect 9255 21184 9271 21248
rect 9335 21184 9351 21248
rect 9415 21184 9423 21248
rect 9103 21183 9423 21184
rect 0 20770 800 20800
rect 1577 20770 1643 20773
rect 0 20768 1643 20770
rect 0 20712 1582 20768
rect 1638 20712 1643 20768
rect 0 20710 1643 20712
rect 0 20680 800 20710
rect 1577 20707 1643 20710
rect 4207 20704 4527 20705
rect 4207 20640 4215 20704
rect 4279 20640 4295 20704
rect 4359 20640 4375 20704
rect 4439 20640 4455 20704
rect 4519 20640 4527 20704
rect 4207 20639 4527 20640
rect 7471 20704 7791 20705
rect 7471 20640 7479 20704
rect 7543 20640 7559 20704
rect 7623 20640 7639 20704
rect 7703 20640 7719 20704
rect 7783 20640 7791 20704
rect 7471 20639 7791 20640
rect 10041 20634 10107 20637
rect 11200 20634 12000 20664
rect 10041 20632 12000 20634
rect 10041 20576 10046 20632
rect 10102 20576 12000 20632
rect 10041 20574 12000 20576
rect 10041 20571 10107 20574
rect 11200 20544 12000 20574
rect 0 20362 800 20392
rect 3509 20362 3575 20365
rect 0 20360 3575 20362
rect 0 20304 3514 20360
rect 3570 20304 3575 20360
rect 0 20302 3575 20304
rect 0 20272 800 20302
rect 3509 20299 3575 20302
rect 2576 20160 2896 20161
rect 2576 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2576 20095 2896 20096
rect 5839 20160 6159 20161
rect 5839 20096 5847 20160
rect 5911 20096 5927 20160
rect 5991 20096 6007 20160
rect 6071 20096 6087 20160
rect 6151 20096 6159 20160
rect 5839 20095 6159 20096
rect 9103 20160 9423 20161
rect 9103 20096 9111 20160
rect 9175 20096 9191 20160
rect 9255 20096 9271 20160
rect 9335 20096 9351 20160
rect 9415 20096 9423 20160
rect 9103 20095 9423 20096
rect 0 19954 800 19984
rect 1669 19954 1735 19957
rect 0 19952 1735 19954
rect 0 19896 1674 19952
rect 1730 19896 1735 19952
rect 0 19894 1735 19896
rect 0 19864 800 19894
rect 1669 19891 1735 19894
rect 4207 19616 4527 19617
rect 0 19546 800 19576
rect 4207 19552 4215 19616
rect 4279 19552 4295 19616
rect 4359 19552 4375 19616
rect 4439 19552 4455 19616
rect 4519 19552 4527 19616
rect 4207 19551 4527 19552
rect 7471 19616 7791 19617
rect 7471 19552 7479 19616
rect 7543 19552 7559 19616
rect 7623 19552 7639 19616
rect 7703 19552 7719 19616
rect 7783 19552 7791 19616
rect 7471 19551 7791 19552
rect 1485 19546 1551 19549
rect 0 19544 1551 19546
rect 0 19488 1490 19544
rect 1546 19488 1551 19544
rect 0 19486 1551 19488
rect 0 19456 800 19486
rect 1485 19483 1551 19486
rect 10041 19410 10107 19413
rect 11200 19410 12000 19440
rect 10041 19408 12000 19410
rect 10041 19352 10046 19408
rect 10102 19352 12000 19408
rect 10041 19350 12000 19352
rect 10041 19347 10107 19350
rect 11200 19320 12000 19350
rect 2576 19072 2896 19073
rect 0 19002 800 19032
rect 2576 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2576 19007 2896 19008
rect 5839 19072 6159 19073
rect 5839 19008 5847 19072
rect 5911 19008 5927 19072
rect 5991 19008 6007 19072
rect 6071 19008 6087 19072
rect 6151 19008 6159 19072
rect 5839 19007 6159 19008
rect 9103 19072 9423 19073
rect 9103 19008 9111 19072
rect 9175 19008 9191 19072
rect 9255 19008 9271 19072
rect 9335 19008 9351 19072
rect 9415 19008 9423 19072
rect 9103 19007 9423 19008
rect 1393 19002 1459 19005
rect 0 19000 1459 19002
rect 0 18944 1398 19000
rect 1454 18944 1459 19000
rect 0 18942 1459 18944
rect 0 18912 800 18942
rect 1393 18939 1459 18942
rect 0 18594 800 18624
rect 3969 18594 4035 18597
rect 0 18592 4035 18594
rect 0 18536 3974 18592
rect 4030 18536 4035 18592
rect 0 18534 4035 18536
rect 0 18504 800 18534
rect 3969 18531 4035 18534
rect 4207 18528 4527 18529
rect 4207 18464 4215 18528
rect 4279 18464 4295 18528
rect 4359 18464 4375 18528
rect 4439 18464 4455 18528
rect 4519 18464 4527 18528
rect 4207 18463 4527 18464
rect 7471 18528 7791 18529
rect 7471 18464 7479 18528
rect 7543 18464 7559 18528
rect 7623 18464 7639 18528
rect 7703 18464 7719 18528
rect 7783 18464 7791 18528
rect 7471 18463 7791 18464
rect 10041 18322 10107 18325
rect 11200 18322 12000 18352
rect 10041 18320 12000 18322
rect 10041 18264 10046 18320
rect 10102 18264 12000 18320
rect 10041 18262 12000 18264
rect 10041 18259 10107 18262
rect 11200 18232 12000 18262
rect 0 18186 800 18216
rect 3509 18186 3575 18189
rect 0 18184 3575 18186
rect 0 18128 3514 18184
rect 3570 18128 3575 18184
rect 0 18126 3575 18128
rect 0 18096 800 18126
rect 3509 18123 3575 18126
rect 2576 17984 2896 17985
rect 2576 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2576 17919 2896 17920
rect 5839 17984 6159 17985
rect 5839 17920 5847 17984
rect 5911 17920 5927 17984
rect 5991 17920 6007 17984
rect 6071 17920 6087 17984
rect 6151 17920 6159 17984
rect 5839 17919 6159 17920
rect 9103 17984 9423 17985
rect 9103 17920 9111 17984
rect 9175 17920 9191 17984
rect 9255 17920 9271 17984
rect 9335 17920 9351 17984
rect 9415 17920 9423 17984
rect 9103 17919 9423 17920
rect 0 17642 800 17672
rect 2865 17642 2931 17645
rect 0 17640 2931 17642
rect 0 17584 2870 17640
rect 2926 17584 2931 17640
rect 0 17582 2931 17584
rect 0 17552 800 17582
rect 2865 17579 2931 17582
rect 4207 17440 4527 17441
rect 4207 17376 4215 17440
rect 4279 17376 4295 17440
rect 4359 17376 4375 17440
rect 4439 17376 4455 17440
rect 4519 17376 4527 17440
rect 4207 17375 4527 17376
rect 7471 17440 7791 17441
rect 7471 17376 7479 17440
rect 7543 17376 7559 17440
rect 7623 17376 7639 17440
rect 7703 17376 7719 17440
rect 7783 17376 7791 17440
rect 7471 17375 7791 17376
rect 1393 17368 1459 17373
rect 1393 17312 1398 17368
rect 1454 17312 1459 17368
rect 1393 17307 1459 17312
rect 0 17234 800 17264
rect 1396 17234 1456 17307
rect 0 17174 1456 17234
rect 10041 17234 10107 17237
rect 11200 17234 12000 17264
rect 10041 17232 12000 17234
rect 10041 17176 10046 17232
rect 10102 17176 12000 17232
rect 10041 17174 12000 17176
rect 0 17144 800 17174
rect 10041 17171 10107 17174
rect 11200 17144 12000 17174
rect 2576 16896 2896 16897
rect 0 16826 800 16856
rect 2576 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2576 16831 2896 16832
rect 5839 16896 6159 16897
rect 5839 16832 5847 16896
rect 5911 16832 5927 16896
rect 5991 16832 6007 16896
rect 6071 16832 6087 16896
rect 6151 16832 6159 16896
rect 5839 16831 6159 16832
rect 9103 16896 9423 16897
rect 9103 16832 9111 16896
rect 9175 16832 9191 16896
rect 9255 16832 9271 16896
rect 9335 16832 9351 16896
rect 9415 16832 9423 16896
rect 9103 16831 9423 16832
rect 933 16826 999 16829
rect 0 16824 999 16826
rect 0 16768 938 16824
rect 994 16768 999 16824
rect 0 16766 999 16768
rect 0 16736 800 16766
rect 933 16763 999 16766
rect 4207 16352 4527 16353
rect 0 16282 800 16312
rect 4207 16288 4215 16352
rect 4279 16288 4295 16352
rect 4359 16288 4375 16352
rect 4439 16288 4455 16352
rect 4519 16288 4527 16352
rect 4207 16287 4527 16288
rect 7471 16352 7791 16353
rect 7471 16288 7479 16352
rect 7543 16288 7559 16352
rect 7623 16288 7639 16352
rect 7703 16288 7719 16352
rect 7783 16288 7791 16352
rect 7471 16287 7791 16288
rect 1393 16282 1459 16285
rect 0 16280 1459 16282
rect 0 16224 1398 16280
rect 1454 16224 1459 16280
rect 0 16222 1459 16224
rect 0 16192 800 16222
rect 1393 16219 1459 16222
rect 10041 16146 10107 16149
rect 11200 16146 12000 16176
rect 10041 16144 12000 16146
rect 10041 16088 10046 16144
rect 10102 16088 12000 16144
rect 10041 16086 12000 16088
rect 10041 16083 10107 16086
rect 11200 16056 12000 16086
rect 0 15874 800 15904
rect 2221 15874 2287 15877
rect 0 15872 2287 15874
rect 0 15816 2226 15872
rect 2282 15816 2287 15872
rect 0 15814 2287 15816
rect 0 15784 800 15814
rect 2221 15811 2287 15814
rect 2576 15808 2896 15809
rect 2576 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2576 15743 2896 15744
rect 5839 15808 6159 15809
rect 5839 15744 5847 15808
rect 5911 15744 5927 15808
rect 5991 15744 6007 15808
rect 6071 15744 6087 15808
rect 6151 15744 6159 15808
rect 5839 15743 6159 15744
rect 9103 15808 9423 15809
rect 9103 15744 9111 15808
rect 9175 15744 9191 15808
rect 9255 15744 9271 15808
rect 9335 15744 9351 15808
rect 9415 15744 9423 15808
rect 9103 15743 9423 15744
rect 0 15466 800 15496
rect 2221 15466 2287 15469
rect 0 15464 2287 15466
rect 0 15408 2226 15464
rect 2282 15408 2287 15464
rect 0 15406 2287 15408
rect 0 15376 800 15406
rect 2221 15403 2287 15406
rect 4207 15264 4527 15265
rect 4207 15200 4215 15264
rect 4279 15200 4295 15264
rect 4359 15200 4375 15264
rect 4439 15200 4455 15264
rect 4519 15200 4527 15264
rect 4207 15199 4527 15200
rect 7471 15264 7791 15265
rect 7471 15200 7479 15264
rect 7543 15200 7559 15264
rect 7623 15200 7639 15264
rect 7703 15200 7719 15264
rect 7783 15200 7791 15264
rect 7471 15199 7791 15200
rect 0 15058 800 15088
rect 1485 15058 1551 15061
rect 0 15056 1551 15058
rect 0 15000 1490 15056
rect 1546 15000 1551 15056
rect 0 14998 1551 15000
rect 0 14968 800 14998
rect 1485 14995 1551 14998
rect 10041 15058 10107 15061
rect 11200 15058 12000 15088
rect 10041 15056 12000 15058
rect 10041 15000 10046 15056
rect 10102 15000 12000 15056
rect 10041 14998 12000 15000
rect 10041 14995 10107 14998
rect 11200 14968 12000 14998
rect 2576 14720 2896 14721
rect 2576 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2576 14655 2896 14656
rect 5839 14720 6159 14721
rect 5839 14656 5847 14720
rect 5911 14656 5927 14720
rect 5991 14656 6007 14720
rect 6071 14656 6087 14720
rect 6151 14656 6159 14720
rect 5839 14655 6159 14656
rect 9103 14720 9423 14721
rect 9103 14656 9111 14720
rect 9175 14656 9191 14720
rect 9255 14656 9271 14720
rect 9335 14656 9351 14720
rect 9415 14656 9423 14720
rect 9103 14655 9423 14656
rect 0 14514 800 14544
rect 1393 14514 1459 14517
rect 0 14512 1459 14514
rect 0 14456 1398 14512
rect 1454 14456 1459 14512
rect 0 14454 1459 14456
rect 0 14424 800 14454
rect 1393 14451 1459 14454
rect 4207 14176 4527 14177
rect 0 14106 800 14136
rect 4207 14112 4215 14176
rect 4279 14112 4295 14176
rect 4359 14112 4375 14176
rect 4439 14112 4455 14176
rect 4519 14112 4527 14176
rect 4207 14111 4527 14112
rect 7471 14176 7791 14177
rect 7471 14112 7479 14176
rect 7543 14112 7559 14176
rect 7623 14112 7639 14176
rect 7703 14112 7719 14176
rect 7783 14112 7791 14176
rect 7471 14111 7791 14112
rect 2313 14106 2379 14109
rect 0 14104 2379 14106
rect 0 14048 2318 14104
rect 2374 14048 2379 14104
rect 0 14046 2379 14048
rect 0 14016 800 14046
rect 2313 14043 2379 14046
rect 10041 13970 10107 13973
rect 11200 13970 12000 14000
rect 10041 13968 12000 13970
rect 10041 13912 10046 13968
rect 10102 13912 12000 13968
rect 10041 13910 12000 13912
rect 10041 13907 10107 13910
rect 11200 13880 12000 13910
rect 0 13698 800 13728
rect 2221 13698 2287 13701
rect 0 13696 2287 13698
rect 0 13640 2226 13696
rect 2282 13640 2287 13696
rect 0 13638 2287 13640
rect 0 13608 800 13638
rect 2221 13635 2287 13638
rect 2576 13632 2896 13633
rect 2576 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2576 13567 2896 13568
rect 5839 13632 6159 13633
rect 5839 13568 5847 13632
rect 5911 13568 5927 13632
rect 5991 13568 6007 13632
rect 6071 13568 6087 13632
rect 6151 13568 6159 13632
rect 5839 13567 6159 13568
rect 9103 13632 9423 13633
rect 9103 13568 9111 13632
rect 9175 13568 9191 13632
rect 9255 13568 9271 13632
rect 9335 13568 9351 13632
rect 9415 13568 9423 13632
rect 9103 13567 9423 13568
rect 0 13154 800 13184
rect 1393 13154 1459 13157
rect 0 13152 1459 13154
rect 0 13096 1398 13152
rect 1454 13096 1459 13152
rect 0 13094 1459 13096
rect 0 13064 800 13094
rect 1393 13091 1459 13094
rect 4207 13088 4527 13089
rect 4207 13024 4215 13088
rect 4279 13024 4295 13088
rect 4359 13024 4375 13088
rect 4439 13024 4455 13088
rect 4519 13024 4527 13088
rect 4207 13023 4527 13024
rect 7471 13088 7791 13089
rect 7471 13024 7479 13088
rect 7543 13024 7559 13088
rect 7623 13024 7639 13088
rect 7703 13024 7719 13088
rect 7783 13024 7791 13088
rect 7471 13023 7791 13024
rect 0 12746 800 12776
rect 2221 12746 2287 12749
rect 0 12744 2287 12746
rect 0 12688 2226 12744
rect 2282 12688 2287 12744
rect 0 12686 2287 12688
rect 0 12656 800 12686
rect 2221 12683 2287 12686
rect 10041 12746 10107 12749
rect 11200 12746 12000 12776
rect 10041 12744 12000 12746
rect 10041 12688 10046 12744
rect 10102 12688 12000 12744
rect 10041 12686 12000 12688
rect 10041 12683 10107 12686
rect 11200 12656 12000 12686
rect 2576 12544 2896 12545
rect 2576 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2576 12479 2896 12480
rect 5839 12544 6159 12545
rect 5839 12480 5847 12544
rect 5911 12480 5927 12544
rect 5991 12480 6007 12544
rect 6071 12480 6087 12544
rect 6151 12480 6159 12544
rect 5839 12479 6159 12480
rect 9103 12544 9423 12545
rect 9103 12480 9111 12544
rect 9175 12480 9191 12544
rect 9255 12480 9271 12544
rect 9335 12480 9351 12544
rect 9415 12480 9423 12544
rect 9103 12479 9423 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 4207 12000 4527 12001
rect 4207 11936 4215 12000
rect 4279 11936 4295 12000
rect 4359 11936 4375 12000
rect 4439 11936 4455 12000
rect 4519 11936 4527 12000
rect 4207 11935 4527 11936
rect 7471 12000 7791 12001
rect 7471 11936 7479 12000
rect 7543 11936 7559 12000
rect 7623 11936 7639 12000
rect 7703 11936 7719 12000
rect 7783 11936 7791 12000
rect 7471 11935 7791 11936
rect 0 11794 800 11824
rect 1393 11794 1459 11797
rect 0 11792 1459 11794
rect 0 11736 1398 11792
rect 1454 11736 1459 11792
rect 0 11734 1459 11736
rect 0 11704 800 11734
rect 1393 11731 1459 11734
rect 10041 11658 10107 11661
rect 11200 11658 12000 11688
rect 10041 11656 12000 11658
rect 10041 11600 10046 11656
rect 10102 11600 12000 11656
rect 10041 11598 12000 11600
rect 10041 11595 10107 11598
rect 11200 11568 12000 11598
rect 2576 11456 2896 11457
rect 0 11386 800 11416
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 11391 2896 11392
rect 5839 11456 6159 11457
rect 5839 11392 5847 11456
rect 5911 11392 5927 11456
rect 5991 11392 6007 11456
rect 6071 11392 6087 11456
rect 6151 11392 6159 11456
rect 5839 11391 6159 11392
rect 9103 11456 9423 11457
rect 9103 11392 9111 11456
rect 9175 11392 9191 11456
rect 9255 11392 9271 11456
rect 9335 11392 9351 11456
rect 9415 11392 9423 11456
rect 9103 11391 9423 11392
rect 1393 11386 1459 11389
rect 0 11384 1459 11386
rect 0 11328 1398 11384
rect 1454 11328 1459 11384
rect 0 11326 1459 11328
rect 0 11296 800 11326
rect 1393 11323 1459 11326
rect 0 10888 800 11008
rect 4207 10912 4527 10913
rect 4207 10848 4215 10912
rect 4279 10848 4295 10912
rect 4359 10848 4375 10912
rect 4439 10848 4455 10912
rect 4519 10848 4527 10912
rect 4207 10847 4527 10848
rect 7471 10912 7791 10913
rect 7471 10848 7479 10912
rect 7543 10848 7559 10912
rect 7623 10848 7639 10912
rect 7703 10848 7719 10912
rect 7783 10848 7791 10912
rect 7471 10847 7791 10848
rect 10041 10570 10107 10573
rect 11200 10570 12000 10600
rect 10041 10568 12000 10570
rect 10041 10512 10046 10568
rect 10102 10512 12000 10568
rect 10041 10510 12000 10512
rect 10041 10507 10107 10510
rect 11200 10480 12000 10510
rect 0 10344 800 10464
rect 2576 10368 2896 10369
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 10303 2896 10304
rect 5839 10368 6159 10369
rect 5839 10304 5847 10368
rect 5911 10304 5927 10368
rect 5991 10304 6007 10368
rect 6071 10304 6087 10368
rect 6151 10304 6159 10368
rect 5839 10303 6159 10304
rect 9103 10368 9423 10369
rect 9103 10304 9111 10368
rect 9175 10304 9191 10368
rect 9255 10304 9271 10368
rect 9335 10304 9351 10368
rect 9415 10304 9423 10368
rect 9103 10303 9423 10304
rect 0 9936 800 10056
rect 4207 9824 4527 9825
rect 4207 9760 4215 9824
rect 4279 9760 4295 9824
rect 4359 9760 4375 9824
rect 4439 9760 4455 9824
rect 4519 9760 4527 9824
rect 4207 9759 4527 9760
rect 7471 9824 7791 9825
rect 7471 9760 7479 9824
rect 7543 9760 7559 9824
rect 7623 9760 7639 9824
rect 7703 9760 7719 9824
rect 7783 9760 7791 9824
rect 7471 9759 7791 9760
rect 0 9528 800 9648
rect 10041 9482 10107 9485
rect 11200 9482 12000 9512
rect 10041 9480 12000 9482
rect 10041 9424 10046 9480
rect 10102 9424 12000 9480
rect 10041 9422 12000 9424
rect 10041 9419 10107 9422
rect 11200 9392 12000 9422
rect 2576 9280 2896 9281
rect 0 9120 800 9240
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 9215 2896 9216
rect 5839 9280 6159 9281
rect 5839 9216 5847 9280
rect 5911 9216 5927 9280
rect 5991 9216 6007 9280
rect 6071 9216 6087 9280
rect 6151 9216 6159 9280
rect 5839 9215 6159 9216
rect 9103 9280 9423 9281
rect 9103 9216 9111 9280
rect 9175 9216 9191 9280
rect 9255 9216 9271 9280
rect 9335 9216 9351 9280
rect 9415 9216 9423 9280
rect 9103 9215 9423 9216
rect 4207 8736 4527 8737
rect 0 8576 800 8696
rect 4207 8672 4215 8736
rect 4279 8672 4295 8736
rect 4359 8672 4375 8736
rect 4439 8672 4455 8736
rect 4519 8672 4527 8736
rect 4207 8671 4527 8672
rect 7471 8736 7791 8737
rect 7471 8672 7479 8736
rect 7543 8672 7559 8736
rect 7623 8672 7639 8736
rect 7703 8672 7719 8736
rect 7783 8672 7791 8736
rect 7471 8671 7791 8672
rect 10041 8394 10107 8397
rect 11200 8394 12000 8424
rect 10041 8392 12000 8394
rect 10041 8336 10046 8392
rect 10102 8336 12000 8392
rect 10041 8334 12000 8336
rect 10041 8331 10107 8334
rect 11200 8304 12000 8334
rect 0 8168 800 8288
rect 2576 8192 2896 8193
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 8127 2896 8128
rect 5839 8192 6159 8193
rect 5839 8128 5847 8192
rect 5911 8128 5927 8192
rect 5991 8128 6007 8192
rect 6071 8128 6087 8192
rect 6151 8128 6159 8192
rect 5839 8127 6159 8128
rect 9103 8192 9423 8193
rect 9103 8128 9111 8192
rect 9175 8128 9191 8192
rect 9255 8128 9271 8192
rect 9335 8128 9351 8192
rect 9415 8128 9423 8192
rect 9103 8127 9423 8128
rect 0 7760 800 7880
rect 4207 7648 4527 7649
rect 4207 7584 4215 7648
rect 4279 7584 4295 7648
rect 4359 7584 4375 7648
rect 4439 7584 4455 7648
rect 4519 7584 4527 7648
rect 4207 7583 4527 7584
rect 7471 7648 7791 7649
rect 7471 7584 7479 7648
rect 7543 7584 7559 7648
rect 7623 7584 7639 7648
rect 7703 7584 7719 7648
rect 7783 7584 7791 7648
rect 7471 7583 7791 7584
rect 0 7216 800 7336
rect 10041 7306 10107 7309
rect 11200 7306 12000 7336
rect 10041 7304 12000 7306
rect 10041 7248 10046 7304
rect 10102 7248 12000 7304
rect 10041 7246 12000 7248
rect 10041 7243 10107 7246
rect 11200 7216 12000 7246
rect 2576 7104 2896 7105
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2576 7039 2896 7040
rect 5839 7104 6159 7105
rect 5839 7040 5847 7104
rect 5911 7040 5927 7104
rect 5991 7040 6007 7104
rect 6071 7040 6087 7104
rect 6151 7040 6159 7104
rect 5839 7039 6159 7040
rect 9103 7104 9423 7105
rect 9103 7040 9111 7104
rect 9175 7040 9191 7104
rect 9255 7040 9271 7104
rect 9335 7040 9351 7104
rect 9415 7040 9423 7104
rect 9103 7039 9423 7040
rect 0 6808 800 6928
rect 4207 6560 4527 6561
rect 0 6400 800 6520
rect 4207 6496 4215 6560
rect 4279 6496 4295 6560
rect 4359 6496 4375 6560
rect 4439 6496 4455 6560
rect 4519 6496 4527 6560
rect 4207 6495 4527 6496
rect 7471 6560 7791 6561
rect 7471 6496 7479 6560
rect 7543 6496 7559 6560
rect 7623 6496 7639 6560
rect 7703 6496 7719 6560
rect 7783 6496 7791 6560
rect 7471 6495 7791 6496
rect 10041 6082 10107 6085
rect 11200 6082 12000 6112
rect 10041 6080 12000 6082
rect 10041 6024 10046 6080
rect 10102 6024 12000 6080
rect 10041 6022 12000 6024
rect 10041 6019 10107 6022
rect 2576 6016 2896 6017
rect 0 5856 800 5976
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 5951 2896 5952
rect 5839 6016 6159 6017
rect 5839 5952 5847 6016
rect 5911 5952 5927 6016
rect 5991 5952 6007 6016
rect 6071 5952 6087 6016
rect 6151 5952 6159 6016
rect 5839 5951 6159 5952
rect 9103 6016 9423 6017
rect 9103 5952 9111 6016
rect 9175 5952 9191 6016
rect 9255 5952 9271 6016
rect 9335 5952 9351 6016
rect 9415 5952 9423 6016
rect 11200 5992 12000 6022
rect 9103 5951 9423 5952
rect 0 5448 800 5568
rect 4207 5472 4527 5473
rect 4207 5408 4215 5472
rect 4279 5408 4295 5472
rect 4359 5408 4375 5472
rect 4439 5408 4455 5472
rect 4519 5408 4527 5472
rect 4207 5407 4527 5408
rect 7471 5472 7791 5473
rect 7471 5408 7479 5472
rect 7543 5408 7559 5472
rect 7623 5408 7639 5472
rect 7703 5408 7719 5472
rect 7783 5408 7791 5472
rect 7471 5407 7791 5408
rect 0 5040 800 5160
rect 10041 4994 10107 4997
rect 11200 4994 12000 5024
rect 10041 4992 12000 4994
rect 10041 4936 10046 4992
rect 10102 4936 12000 4992
rect 10041 4934 12000 4936
rect 10041 4931 10107 4934
rect 2576 4928 2896 4929
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 4863 2896 4864
rect 5839 4928 6159 4929
rect 5839 4864 5847 4928
rect 5911 4864 5927 4928
rect 5991 4864 6007 4928
rect 6071 4864 6087 4928
rect 6151 4864 6159 4928
rect 5839 4863 6159 4864
rect 9103 4928 9423 4929
rect 9103 4864 9111 4928
rect 9175 4864 9191 4928
rect 9255 4864 9271 4928
rect 9335 4864 9351 4928
rect 9415 4864 9423 4928
rect 11200 4904 12000 4934
rect 9103 4863 9423 4864
rect 0 4632 800 4752
rect 4207 4384 4527 4385
rect 4207 4320 4215 4384
rect 4279 4320 4295 4384
rect 4359 4320 4375 4384
rect 4439 4320 4455 4384
rect 4519 4320 4527 4384
rect 4207 4319 4527 4320
rect 7471 4384 7791 4385
rect 7471 4320 7479 4384
rect 7543 4320 7559 4384
rect 7623 4320 7639 4384
rect 7703 4320 7719 4384
rect 7783 4320 7791 4384
rect 7471 4319 7791 4320
rect 0 4088 800 4208
rect 10041 3906 10107 3909
rect 11200 3906 12000 3936
rect 10041 3904 12000 3906
rect 10041 3848 10046 3904
rect 10102 3848 12000 3904
rect 10041 3846 12000 3848
rect 10041 3843 10107 3846
rect 2576 3840 2896 3841
rect 0 3770 800 3800
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 3775 2896 3776
rect 5839 3840 6159 3841
rect 5839 3776 5847 3840
rect 5911 3776 5927 3840
rect 5991 3776 6007 3840
rect 6071 3776 6087 3840
rect 6151 3776 6159 3840
rect 5839 3775 6159 3776
rect 9103 3840 9423 3841
rect 9103 3776 9111 3840
rect 9175 3776 9191 3840
rect 9255 3776 9271 3840
rect 9335 3776 9351 3840
rect 9415 3776 9423 3840
rect 11200 3816 12000 3846
rect 9103 3775 9423 3776
rect 1393 3770 1459 3773
rect 0 3768 1459 3770
rect 0 3712 1398 3768
rect 1454 3712 1459 3768
rect 0 3710 1459 3712
rect 0 3680 800 3710
rect 1393 3707 1459 3710
rect 0 3362 800 3392
rect 1209 3362 1275 3365
rect 0 3360 1275 3362
rect 0 3304 1214 3360
rect 1270 3304 1275 3360
rect 0 3302 1275 3304
rect 0 3272 800 3302
rect 1209 3299 1275 3302
rect 4207 3296 4527 3297
rect 4207 3232 4215 3296
rect 4279 3232 4295 3296
rect 4359 3232 4375 3296
rect 4439 3232 4455 3296
rect 4519 3232 4527 3296
rect 4207 3231 4527 3232
rect 7471 3296 7791 3297
rect 7471 3232 7479 3296
rect 7543 3232 7559 3296
rect 7623 3232 7639 3296
rect 7703 3232 7719 3296
rect 7783 3232 7791 3296
rect 7471 3231 7791 3232
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 10041 2818 10107 2821
rect 11200 2818 12000 2848
rect 10041 2816 12000 2818
rect 10041 2760 10046 2816
rect 10102 2760 12000 2816
rect 10041 2758 12000 2760
rect 10041 2755 10107 2758
rect 2576 2752 2896 2753
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2687 2896 2688
rect 5839 2752 6159 2753
rect 5839 2688 5847 2752
rect 5911 2688 5927 2752
rect 5991 2688 6007 2752
rect 6071 2688 6087 2752
rect 6151 2688 6159 2752
rect 5839 2687 6159 2688
rect 9103 2752 9423 2753
rect 9103 2688 9111 2752
rect 9175 2688 9191 2752
rect 9255 2688 9271 2752
rect 9335 2688 9351 2752
rect 9415 2688 9423 2752
rect 11200 2728 12000 2758
rect 9103 2687 9423 2688
rect 0 2410 800 2440
rect 1393 2410 1459 2413
rect 0 2408 1459 2410
rect 0 2352 1398 2408
rect 1454 2352 1459 2408
rect 0 2350 1459 2352
rect 0 2320 800 2350
rect 1393 2347 1459 2350
rect 4207 2208 4527 2209
rect 4207 2144 4215 2208
rect 4279 2144 4295 2208
rect 4359 2144 4375 2208
rect 4439 2144 4455 2208
rect 4519 2144 4527 2208
rect 4207 2143 4527 2144
rect 7471 2208 7791 2209
rect 7471 2144 7479 2208
rect 7543 2144 7559 2208
rect 7623 2144 7639 2208
rect 7703 2144 7719 2208
rect 7783 2144 7791 2208
rect 7471 2143 7791 2144
rect 0 2002 800 2032
rect 2773 2002 2839 2005
rect 0 2000 2839 2002
rect 0 1944 2778 2000
rect 2834 1944 2839 2000
rect 0 1942 2839 1944
rect 0 1912 800 1942
rect 2773 1939 2839 1942
rect 10041 1730 10107 1733
rect 11200 1730 12000 1760
rect 10041 1728 12000 1730
rect 10041 1672 10046 1728
rect 10102 1672 12000 1728
rect 10041 1670 12000 1672
rect 10041 1667 10107 1670
rect 11200 1640 12000 1670
rect 0 1458 800 1488
rect 1301 1458 1367 1461
rect 0 1456 1367 1458
rect 0 1400 1306 1456
rect 1362 1400 1367 1456
rect 0 1398 1367 1400
rect 0 1368 800 1398
rect 1301 1395 1367 1398
rect 0 1050 800 1080
rect 2037 1050 2103 1053
rect 0 1048 2103 1050
rect 0 992 2042 1048
rect 2098 992 2103 1048
rect 0 990 2103 992
rect 0 960 800 990
rect 2037 987 2103 990
rect 0 552 800 672
rect 10961 642 11027 645
rect 11200 642 12000 672
rect 10961 640 12000 642
rect 10961 584 10966 640
rect 11022 584 12000 640
rect 10961 582 12000 584
rect 10961 579 11027 582
rect 11200 552 12000 582
rect 0 144 800 264
<< via3 >>
rect 2584 77820 2648 77824
rect 2584 77764 2588 77820
rect 2588 77764 2644 77820
rect 2644 77764 2648 77820
rect 2584 77760 2648 77764
rect 2664 77820 2728 77824
rect 2664 77764 2668 77820
rect 2668 77764 2724 77820
rect 2724 77764 2728 77820
rect 2664 77760 2728 77764
rect 2744 77820 2808 77824
rect 2744 77764 2748 77820
rect 2748 77764 2804 77820
rect 2804 77764 2808 77820
rect 2744 77760 2808 77764
rect 2824 77820 2888 77824
rect 2824 77764 2828 77820
rect 2828 77764 2884 77820
rect 2884 77764 2888 77820
rect 2824 77760 2888 77764
rect 5847 77820 5911 77824
rect 5847 77764 5851 77820
rect 5851 77764 5907 77820
rect 5907 77764 5911 77820
rect 5847 77760 5911 77764
rect 5927 77820 5991 77824
rect 5927 77764 5931 77820
rect 5931 77764 5987 77820
rect 5987 77764 5991 77820
rect 5927 77760 5991 77764
rect 6007 77820 6071 77824
rect 6007 77764 6011 77820
rect 6011 77764 6067 77820
rect 6067 77764 6071 77820
rect 6007 77760 6071 77764
rect 6087 77820 6151 77824
rect 6087 77764 6091 77820
rect 6091 77764 6147 77820
rect 6147 77764 6151 77820
rect 6087 77760 6151 77764
rect 9111 77820 9175 77824
rect 9111 77764 9115 77820
rect 9115 77764 9171 77820
rect 9171 77764 9175 77820
rect 9111 77760 9175 77764
rect 9191 77820 9255 77824
rect 9191 77764 9195 77820
rect 9195 77764 9251 77820
rect 9251 77764 9255 77820
rect 9191 77760 9255 77764
rect 9271 77820 9335 77824
rect 9271 77764 9275 77820
rect 9275 77764 9331 77820
rect 9331 77764 9335 77820
rect 9271 77760 9335 77764
rect 9351 77820 9415 77824
rect 9351 77764 9355 77820
rect 9355 77764 9411 77820
rect 9411 77764 9415 77820
rect 9351 77760 9415 77764
rect 4215 77276 4279 77280
rect 4215 77220 4219 77276
rect 4219 77220 4275 77276
rect 4275 77220 4279 77276
rect 4215 77216 4279 77220
rect 4295 77276 4359 77280
rect 4295 77220 4299 77276
rect 4299 77220 4355 77276
rect 4355 77220 4359 77276
rect 4295 77216 4359 77220
rect 4375 77276 4439 77280
rect 4375 77220 4379 77276
rect 4379 77220 4435 77276
rect 4435 77220 4439 77276
rect 4375 77216 4439 77220
rect 4455 77276 4519 77280
rect 4455 77220 4459 77276
rect 4459 77220 4515 77276
rect 4515 77220 4519 77276
rect 4455 77216 4519 77220
rect 7479 77276 7543 77280
rect 7479 77220 7483 77276
rect 7483 77220 7539 77276
rect 7539 77220 7543 77276
rect 7479 77216 7543 77220
rect 7559 77276 7623 77280
rect 7559 77220 7563 77276
rect 7563 77220 7619 77276
rect 7619 77220 7623 77276
rect 7559 77216 7623 77220
rect 7639 77276 7703 77280
rect 7639 77220 7643 77276
rect 7643 77220 7699 77276
rect 7699 77220 7703 77276
rect 7639 77216 7703 77220
rect 7719 77276 7783 77280
rect 7719 77220 7723 77276
rect 7723 77220 7779 77276
rect 7779 77220 7783 77276
rect 7719 77216 7783 77220
rect 2584 76732 2648 76736
rect 2584 76676 2588 76732
rect 2588 76676 2644 76732
rect 2644 76676 2648 76732
rect 2584 76672 2648 76676
rect 2664 76732 2728 76736
rect 2664 76676 2668 76732
rect 2668 76676 2724 76732
rect 2724 76676 2728 76732
rect 2664 76672 2728 76676
rect 2744 76732 2808 76736
rect 2744 76676 2748 76732
rect 2748 76676 2804 76732
rect 2804 76676 2808 76732
rect 2744 76672 2808 76676
rect 2824 76732 2888 76736
rect 2824 76676 2828 76732
rect 2828 76676 2884 76732
rect 2884 76676 2888 76732
rect 2824 76672 2888 76676
rect 5847 76732 5911 76736
rect 5847 76676 5851 76732
rect 5851 76676 5907 76732
rect 5907 76676 5911 76732
rect 5847 76672 5911 76676
rect 5927 76732 5991 76736
rect 5927 76676 5931 76732
rect 5931 76676 5987 76732
rect 5987 76676 5991 76732
rect 5927 76672 5991 76676
rect 6007 76732 6071 76736
rect 6007 76676 6011 76732
rect 6011 76676 6067 76732
rect 6067 76676 6071 76732
rect 6007 76672 6071 76676
rect 6087 76732 6151 76736
rect 6087 76676 6091 76732
rect 6091 76676 6147 76732
rect 6147 76676 6151 76732
rect 6087 76672 6151 76676
rect 9111 76732 9175 76736
rect 9111 76676 9115 76732
rect 9115 76676 9171 76732
rect 9171 76676 9175 76732
rect 9111 76672 9175 76676
rect 9191 76732 9255 76736
rect 9191 76676 9195 76732
rect 9195 76676 9251 76732
rect 9251 76676 9255 76732
rect 9191 76672 9255 76676
rect 9271 76732 9335 76736
rect 9271 76676 9275 76732
rect 9275 76676 9331 76732
rect 9331 76676 9335 76732
rect 9271 76672 9335 76676
rect 9351 76732 9415 76736
rect 9351 76676 9355 76732
rect 9355 76676 9411 76732
rect 9411 76676 9415 76732
rect 9351 76672 9415 76676
rect 4215 76188 4279 76192
rect 4215 76132 4219 76188
rect 4219 76132 4275 76188
rect 4275 76132 4279 76188
rect 4215 76128 4279 76132
rect 4295 76188 4359 76192
rect 4295 76132 4299 76188
rect 4299 76132 4355 76188
rect 4355 76132 4359 76188
rect 4295 76128 4359 76132
rect 4375 76188 4439 76192
rect 4375 76132 4379 76188
rect 4379 76132 4435 76188
rect 4435 76132 4439 76188
rect 4375 76128 4439 76132
rect 4455 76188 4519 76192
rect 4455 76132 4459 76188
rect 4459 76132 4515 76188
rect 4515 76132 4519 76188
rect 4455 76128 4519 76132
rect 7479 76188 7543 76192
rect 7479 76132 7483 76188
rect 7483 76132 7539 76188
rect 7539 76132 7543 76188
rect 7479 76128 7543 76132
rect 7559 76188 7623 76192
rect 7559 76132 7563 76188
rect 7563 76132 7619 76188
rect 7619 76132 7623 76188
rect 7559 76128 7623 76132
rect 7639 76188 7703 76192
rect 7639 76132 7643 76188
rect 7643 76132 7699 76188
rect 7699 76132 7703 76188
rect 7639 76128 7703 76132
rect 7719 76188 7783 76192
rect 7719 76132 7723 76188
rect 7723 76132 7779 76188
rect 7779 76132 7783 76188
rect 7719 76128 7783 76132
rect 2584 75644 2648 75648
rect 2584 75588 2588 75644
rect 2588 75588 2644 75644
rect 2644 75588 2648 75644
rect 2584 75584 2648 75588
rect 2664 75644 2728 75648
rect 2664 75588 2668 75644
rect 2668 75588 2724 75644
rect 2724 75588 2728 75644
rect 2664 75584 2728 75588
rect 2744 75644 2808 75648
rect 2744 75588 2748 75644
rect 2748 75588 2804 75644
rect 2804 75588 2808 75644
rect 2744 75584 2808 75588
rect 2824 75644 2888 75648
rect 2824 75588 2828 75644
rect 2828 75588 2884 75644
rect 2884 75588 2888 75644
rect 2824 75584 2888 75588
rect 5847 75644 5911 75648
rect 5847 75588 5851 75644
rect 5851 75588 5907 75644
rect 5907 75588 5911 75644
rect 5847 75584 5911 75588
rect 5927 75644 5991 75648
rect 5927 75588 5931 75644
rect 5931 75588 5987 75644
rect 5987 75588 5991 75644
rect 5927 75584 5991 75588
rect 6007 75644 6071 75648
rect 6007 75588 6011 75644
rect 6011 75588 6067 75644
rect 6067 75588 6071 75644
rect 6007 75584 6071 75588
rect 6087 75644 6151 75648
rect 6087 75588 6091 75644
rect 6091 75588 6147 75644
rect 6147 75588 6151 75644
rect 6087 75584 6151 75588
rect 9111 75644 9175 75648
rect 9111 75588 9115 75644
rect 9115 75588 9171 75644
rect 9171 75588 9175 75644
rect 9111 75584 9175 75588
rect 9191 75644 9255 75648
rect 9191 75588 9195 75644
rect 9195 75588 9251 75644
rect 9251 75588 9255 75644
rect 9191 75584 9255 75588
rect 9271 75644 9335 75648
rect 9271 75588 9275 75644
rect 9275 75588 9331 75644
rect 9331 75588 9335 75644
rect 9271 75584 9335 75588
rect 9351 75644 9415 75648
rect 9351 75588 9355 75644
rect 9355 75588 9411 75644
rect 9411 75588 9415 75644
rect 9351 75584 9415 75588
rect 4215 75100 4279 75104
rect 4215 75044 4219 75100
rect 4219 75044 4275 75100
rect 4275 75044 4279 75100
rect 4215 75040 4279 75044
rect 4295 75100 4359 75104
rect 4295 75044 4299 75100
rect 4299 75044 4355 75100
rect 4355 75044 4359 75100
rect 4295 75040 4359 75044
rect 4375 75100 4439 75104
rect 4375 75044 4379 75100
rect 4379 75044 4435 75100
rect 4435 75044 4439 75100
rect 4375 75040 4439 75044
rect 4455 75100 4519 75104
rect 4455 75044 4459 75100
rect 4459 75044 4515 75100
rect 4515 75044 4519 75100
rect 4455 75040 4519 75044
rect 7479 75100 7543 75104
rect 7479 75044 7483 75100
rect 7483 75044 7539 75100
rect 7539 75044 7543 75100
rect 7479 75040 7543 75044
rect 7559 75100 7623 75104
rect 7559 75044 7563 75100
rect 7563 75044 7619 75100
rect 7619 75044 7623 75100
rect 7559 75040 7623 75044
rect 7639 75100 7703 75104
rect 7639 75044 7643 75100
rect 7643 75044 7699 75100
rect 7699 75044 7703 75100
rect 7639 75040 7703 75044
rect 7719 75100 7783 75104
rect 7719 75044 7723 75100
rect 7723 75044 7779 75100
rect 7779 75044 7783 75100
rect 7719 75040 7783 75044
rect 2584 74556 2648 74560
rect 2584 74500 2588 74556
rect 2588 74500 2644 74556
rect 2644 74500 2648 74556
rect 2584 74496 2648 74500
rect 2664 74556 2728 74560
rect 2664 74500 2668 74556
rect 2668 74500 2724 74556
rect 2724 74500 2728 74556
rect 2664 74496 2728 74500
rect 2744 74556 2808 74560
rect 2744 74500 2748 74556
rect 2748 74500 2804 74556
rect 2804 74500 2808 74556
rect 2744 74496 2808 74500
rect 2824 74556 2888 74560
rect 2824 74500 2828 74556
rect 2828 74500 2884 74556
rect 2884 74500 2888 74556
rect 2824 74496 2888 74500
rect 5847 74556 5911 74560
rect 5847 74500 5851 74556
rect 5851 74500 5907 74556
rect 5907 74500 5911 74556
rect 5847 74496 5911 74500
rect 5927 74556 5991 74560
rect 5927 74500 5931 74556
rect 5931 74500 5987 74556
rect 5987 74500 5991 74556
rect 5927 74496 5991 74500
rect 6007 74556 6071 74560
rect 6007 74500 6011 74556
rect 6011 74500 6067 74556
rect 6067 74500 6071 74556
rect 6007 74496 6071 74500
rect 6087 74556 6151 74560
rect 6087 74500 6091 74556
rect 6091 74500 6147 74556
rect 6147 74500 6151 74556
rect 6087 74496 6151 74500
rect 9111 74556 9175 74560
rect 9111 74500 9115 74556
rect 9115 74500 9171 74556
rect 9171 74500 9175 74556
rect 9111 74496 9175 74500
rect 9191 74556 9255 74560
rect 9191 74500 9195 74556
rect 9195 74500 9251 74556
rect 9251 74500 9255 74556
rect 9191 74496 9255 74500
rect 9271 74556 9335 74560
rect 9271 74500 9275 74556
rect 9275 74500 9331 74556
rect 9331 74500 9335 74556
rect 9271 74496 9335 74500
rect 9351 74556 9415 74560
rect 9351 74500 9355 74556
rect 9355 74500 9411 74556
rect 9411 74500 9415 74556
rect 9351 74496 9415 74500
rect 4215 74012 4279 74016
rect 4215 73956 4219 74012
rect 4219 73956 4275 74012
rect 4275 73956 4279 74012
rect 4215 73952 4279 73956
rect 4295 74012 4359 74016
rect 4295 73956 4299 74012
rect 4299 73956 4355 74012
rect 4355 73956 4359 74012
rect 4295 73952 4359 73956
rect 4375 74012 4439 74016
rect 4375 73956 4379 74012
rect 4379 73956 4435 74012
rect 4435 73956 4439 74012
rect 4375 73952 4439 73956
rect 4455 74012 4519 74016
rect 4455 73956 4459 74012
rect 4459 73956 4515 74012
rect 4515 73956 4519 74012
rect 4455 73952 4519 73956
rect 7479 74012 7543 74016
rect 7479 73956 7483 74012
rect 7483 73956 7539 74012
rect 7539 73956 7543 74012
rect 7479 73952 7543 73956
rect 7559 74012 7623 74016
rect 7559 73956 7563 74012
rect 7563 73956 7619 74012
rect 7619 73956 7623 74012
rect 7559 73952 7623 73956
rect 7639 74012 7703 74016
rect 7639 73956 7643 74012
rect 7643 73956 7699 74012
rect 7699 73956 7703 74012
rect 7639 73952 7703 73956
rect 7719 74012 7783 74016
rect 7719 73956 7723 74012
rect 7723 73956 7779 74012
rect 7779 73956 7783 74012
rect 7719 73952 7783 73956
rect 2584 73468 2648 73472
rect 2584 73412 2588 73468
rect 2588 73412 2644 73468
rect 2644 73412 2648 73468
rect 2584 73408 2648 73412
rect 2664 73468 2728 73472
rect 2664 73412 2668 73468
rect 2668 73412 2724 73468
rect 2724 73412 2728 73468
rect 2664 73408 2728 73412
rect 2744 73468 2808 73472
rect 2744 73412 2748 73468
rect 2748 73412 2804 73468
rect 2804 73412 2808 73468
rect 2744 73408 2808 73412
rect 2824 73468 2888 73472
rect 2824 73412 2828 73468
rect 2828 73412 2884 73468
rect 2884 73412 2888 73468
rect 2824 73408 2888 73412
rect 5847 73468 5911 73472
rect 5847 73412 5851 73468
rect 5851 73412 5907 73468
rect 5907 73412 5911 73468
rect 5847 73408 5911 73412
rect 5927 73468 5991 73472
rect 5927 73412 5931 73468
rect 5931 73412 5987 73468
rect 5987 73412 5991 73468
rect 5927 73408 5991 73412
rect 6007 73468 6071 73472
rect 6007 73412 6011 73468
rect 6011 73412 6067 73468
rect 6067 73412 6071 73468
rect 6007 73408 6071 73412
rect 6087 73468 6151 73472
rect 6087 73412 6091 73468
rect 6091 73412 6147 73468
rect 6147 73412 6151 73468
rect 6087 73408 6151 73412
rect 9111 73468 9175 73472
rect 9111 73412 9115 73468
rect 9115 73412 9171 73468
rect 9171 73412 9175 73468
rect 9111 73408 9175 73412
rect 9191 73468 9255 73472
rect 9191 73412 9195 73468
rect 9195 73412 9251 73468
rect 9251 73412 9255 73468
rect 9191 73408 9255 73412
rect 9271 73468 9335 73472
rect 9271 73412 9275 73468
rect 9275 73412 9331 73468
rect 9331 73412 9335 73468
rect 9271 73408 9335 73412
rect 9351 73468 9415 73472
rect 9351 73412 9355 73468
rect 9355 73412 9411 73468
rect 9411 73412 9415 73468
rect 9351 73408 9415 73412
rect 4215 72924 4279 72928
rect 4215 72868 4219 72924
rect 4219 72868 4275 72924
rect 4275 72868 4279 72924
rect 4215 72864 4279 72868
rect 4295 72924 4359 72928
rect 4295 72868 4299 72924
rect 4299 72868 4355 72924
rect 4355 72868 4359 72924
rect 4295 72864 4359 72868
rect 4375 72924 4439 72928
rect 4375 72868 4379 72924
rect 4379 72868 4435 72924
rect 4435 72868 4439 72924
rect 4375 72864 4439 72868
rect 4455 72924 4519 72928
rect 4455 72868 4459 72924
rect 4459 72868 4515 72924
rect 4515 72868 4519 72924
rect 4455 72864 4519 72868
rect 7479 72924 7543 72928
rect 7479 72868 7483 72924
rect 7483 72868 7539 72924
rect 7539 72868 7543 72924
rect 7479 72864 7543 72868
rect 7559 72924 7623 72928
rect 7559 72868 7563 72924
rect 7563 72868 7619 72924
rect 7619 72868 7623 72924
rect 7559 72864 7623 72868
rect 7639 72924 7703 72928
rect 7639 72868 7643 72924
rect 7643 72868 7699 72924
rect 7699 72868 7703 72924
rect 7639 72864 7703 72868
rect 7719 72924 7783 72928
rect 7719 72868 7723 72924
rect 7723 72868 7779 72924
rect 7779 72868 7783 72924
rect 7719 72864 7783 72868
rect 2584 72380 2648 72384
rect 2584 72324 2588 72380
rect 2588 72324 2644 72380
rect 2644 72324 2648 72380
rect 2584 72320 2648 72324
rect 2664 72380 2728 72384
rect 2664 72324 2668 72380
rect 2668 72324 2724 72380
rect 2724 72324 2728 72380
rect 2664 72320 2728 72324
rect 2744 72380 2808 72384
rect 2744 72324 2748 72380
rect 2748 72324 2804 72380
rect 2804 72324 2808 72380
rect 2744 72320 2808 72324
rect 2824 72380 2888 72384
rect 2824 72324 2828 72380
rect 2828 72324 2884 72380
rect 2884 72324 2888 72380
rect 2824 72320 2888 72324
rect 5847 72380 5911 72384
rect 5847 72324 5851 72380
rect 5851 72324 5907 72380
rect 5907 72324 5911 72380
rect 5847 72320 5911 72324
rect 5927 72380 5991 72384
rect 5927 72324 5931 72380
rect 5931 72324 5987 72380
rect 5987 72324 5991 72380
rect 5927 72320 5991 72324
rect 6007 72380 6071 72384
rect 6007 72324 6011 72380
rect 6011 72324 6067 72380
rect 6067 72324 6071 72380
rect 6007 72320 6071 72324
rect 6087 72380 6151 72384
rect 6087 72324 6091 72380
rect 6091 72324 6147 72380
rect 6147 72324 6151 72380
rect 6087 72320 6151 72324
rect 9111 72380 9175 72384
rect 9111 72324 9115 72380
rect 9115 72324 9171 72380
rect 9171 72324 9175 72380
rect 9111 72320 9175 72324
rect 9191 72380 9255 72384
rect 9191 72324 9195 72380
rect 9195 72324 9251 72380
rect 9251 72324 9255 72380
rect 9191 72320 9255 72324
rect 9271 72380 9335 72384
rect 9271 72324 9275 72380
rect 9275 72324 9331 72380
rect 9331 72324 9335 72380
rect 9271 72320 9335 72324
rect 9351 72380 9415 72384
rect 9351 72324 9355 72380
rect 9355 72324 9411 72380
rect 9411 72324 9415 72380
rect 9351 72320 9415 72324
rect 4215 71836 4279 71840
rect 4215 71780 4219 71836
rect 4219 71780 4275 71836
rect 4275 71780 4279 71836
rect 4215 71776 4279 71780
rect 4295 71836 4359 71840
rect 4295 71780 4299 71836
rect 4299 71780 4355 71836
rect 4355 71780 4359 71836
rect 4295 71776 4359 71780
rect 4375 71836 4439 71840
rect 4375 71780 4379 71836
rect 4379 71780 4435 71836
rect 4435 71780 4439 71836
rect 4375 71776 4439 71780
rect 4455 71836 4519 71840
rect 4455 71780 4459 71836
rect 4459 71780 4515 71836
rect 4515 71780 4519 71836
rect 4455 71776 4519 71780
rect 7479 71836 7543 71840
rect 7479 71780 7483 71836
rect 7483 71780 7539 71836
rect 7539 71780 7543 71836
rect 7479 71776 7543 71780
rect 7559 71836 7623 71840
rect 7559 71780 7563 71836
rect 7563 71780 7619 71836
rect 7619 71780 7623 71836
rect 7559 71776 7623 71780
rect 7639 71836 7703 71840
rect 7639 71780 7643 71836
rect 7643 71780 7699 71836
rect 7699 71780 7703 71836
rect 7639 71776 7703 71780
rect 7719 71836 7783 71840
rect 7719 71780 7723 71836
rect 7723 71780 7779 71836
rect 7779 71780 7783 71836
rect 7719 71776 7783 71780
rect 2584 71292 2648 71296
rect 2584 71236 2588 71292
rect 2588 71236 2644 71292
rect 2644 71236 2648 71292
rect 2584 71232 2648 71236
rect 2664 71292 2728 71296
rect 2664 71236 2668 71292
rect 2668 71236 2724 71292
rect 2724 71236 2728 71292
rect 2664 71232 2728 71236
rect 2744 71292 2808 71296
rect 2744 71236 2748 71292
rect 2748 71236 2804 71292
rect 2804 71236 2808 71292
rect 2744 71232 2808 71236
rect 2824 71292 2888 71296
rect 2824 71236 2828 71292
rect 2828 71236 2884 71292
rect 2884 71236 2888 71292
rect 2824 71232 2888 71236
rect 5847 71292 5911 71296
rect 5847 71236 5851 71292
rect 5851 71236 5907 71292
rect 5907 71236 5911 71292
rect 5847 71232 5911 71236
rect 5927 71292 5991 71296
rect 5927 71236 5931 71292
rect 5931 71236 5987 71292
rect 5987 71236 5991 71292
rect 5927 71232 5991 71236
rect 6007 71292 6071 71296
rect 6007 71236 6011 71292
rect 6011 71236 6067 71292
rect 6067 71236 6071 71292
rect 6007 71232 6071 71236
rect 6087 71292 6151 71296
rect 6087 71236 6091 71292
rect 6091 71236 6147 71292
rect 6147 71236 6151 71292
rect 6087 71232 6151 71236
rect 9111 71292 9175 71296
rect 9111 71236 9115 71292
rect 9115 71236 9171 71292
rect 9171 71236 9175 71292
rect 9111 71232 9175 71236
rect 9191 71292 9255 71296
rect 9191 71236 9195 71292
rect 9195 71236 9251 71292
rect 9251 71236 9255 71292
rect 9191 71232 9255 71236
rect 9271 71292 9335 71296
rect 9271 71236 9275 71292
rect 9275 71236 9331 71292
rect 9331 71236 9335 71292
rect 9271 71232 9335 71236
rect 9351 71292 9415 71296
rect 9351 71236 9355 71292
rect 9355 71236 9411 71292
rect 9411 71236 9415 71292
rect 9351 71232 9415 71236
rect 4215 70748 4279 70752
rect 4215 70692 4219 70748
rect 4219 70692 4275 70748
rect 4275 70692 4279 70748
rect 4215 70688 4279 70692
rect 4295 70748 4359 70752
rect 4295 70692 4299 70748
rect 4299 70692 4355 70748
rect 4355 70692 4359 70748
rect 4295 70688 4359 70692
rect 4375 70748 4439 70752
rect 4375 70692 4379 70748
rect 4379 70692 4435 70748
rect 4435 70692 4439 70748
rect 4375 70688 4439 70692
rect 4455 70748 4519 70752
rect 4455 70692 4459 70748
rect 4459 70692 4515 70748
rect 4515 70692 4519 70748
rect 4455 70688 4519 70692
rect 7479 70748 7543 70752
rect 7479 70692 7483 70748
rect 7483 70692 7539 70748
rect 7539 70692 7543 70748
rect 7479 70688 7543 70692
rect 7559 70748 7623 70752
rect 7559 70692 7563 70748
rect 7563 70692 7619 70748
rect 7619 70692 7623 70748
rect 7559 70688 7623 70692
rect 7639 70748 7703 70752
rect 7639 70692 7643 70748
rect 7643 70692 7699 70748
rect 7699 70692 7703 70748
rect 7639 70688 7703 70692
rect 7719 70748 7783 70752
rect 7719 70692 7723 70748
rect 7723 70692 7779 70748
rect 7779 70692 7783 70748
rect 7719 70688 7783 70692
rect 1532 70484 1596 70548
rect 2584 70204 2648 70208
rect 2584 70148 2588 70204
rect 2588 70148 2644 70204
rect 2644 70148 2648 70204
rect 2584 70144 2648 70148
rect 2664 70204 2728 70208
rect 2664 70148 2668 70204
rect 2668 70148 2724 70204
rect 2724 70148 2728 70204
rect 2664 70144 2728 70148
rect 2744 70204 2808 70208
rect 2744 70148 2748 70204
rect 2748 70148 2804 70204
rect 2804 70148 2808 70204
rect 2744 70144 2808 70148
rect 2824 70204 2888 70208
rect 2824 70148 2828 70204
rect 2828 70148 2884 70204
rect 2884 70148 2888 70204
rect 2824 70144 2888 70148
rect 5847 70204 5911 70208
rect 5847 70148 5851 70204
rect 5851 70148 5907 70204
rect 5907 70148 5911 70204
rect 5847 70144 5911 70148
rect 5927 70204 5991 70208
rect 5927 70148 5931 70204
rect 5931 70148 5987 70204
rect 5987 70148 5991 70204
rect 5927 70144 5991 70148
rect 6007 70204 6071 70208
rect 6007 70148 6011 70204
rect 6011 70148 6067 70204
rect 6067 70148 6071 70204
rect 6007 70144 6071 70148
rect 6087 70204 6151 70208
rect 6087 70148 6091 70204
rect 6091 70148 6147 70204
rect 6147 70148 6151 70204
rect 6087 70144 6151 70148
rect 9111 70204 9175 70208
rect 9111 70148 9115 70204
rect 9115 70148 9171 70204
rect 9171 70148 9175 70204
rect 9111 70144 9175 70148
rect 9191 70204 9255 70208
rect 9191 70148 9195 70204
rect 9195 70148 9251 70204
rect 9251 70148 9255 70204
rect 9191 70144 9255 70148
rect 9271 70204 9335 70208
rect 9271 70148 9275 70204
rect 9275 70148 9331 70204
rect 9331 70148 9335 70204
rect 9271 70144 9335 70148
rect 9351 70204 9415 70208
rect 9351 70148 9355 70204
rect 9355 70148 9411 70204
rect 9411 70148 9415 70204
rect 9351 70144 9415 70148
rect 4215 69660 4279 69664
rect 4215 69604 4219 69660
rect 4219 69604 4275 69660
rect 4275 69604 4279 69660
rect 4215 69600 4279 69604
rect 4295 69660 4359 69664
rect 4295 69604 4299 69660
rect 4299 69604 4355 69660
rect 4355 69604 4359 69660
rect 4295 69600 4359 69604
rect 4375 69660 4439 69664
rect 4375 69604 4379 69660
rect 4379 69604 4435 69660
rect 4435 69604 4439 69660
rect 4375 69600 4439 69604
rect 4455 69660 4519 69664
rect 4455 69604 4459 69660
rect 4459 69604 4515 69660
rect 4515 69604 4519 69660
rect 4455 69600 4519 69604
rect 7479 69660 7543 69664
rect 7479 69604 7483 69660
rect 7483 69604 7539 69660
rect 7539 69604 7543 69660
rect 7479 69600 7543 69604
rect 7559 69660 7623 69664
rect 7559 69604 7563 69660
rect 7563 69604 7619 69660
rect 7619 69604 7623 69660
rect 7559 69600 7623 69604
rect 7639 69660 7703 69664
rect 7639 69604 7643 69660
rect 7643 69604 7699 69660
rect 7699 69604 7703 69660
rect 7639 69600 7703 69604
rect 7719 69660 7783 69664
rect 7719 69604 7723 69660
rect 7723 69604 7779 69660
rect 7779 69604 7783 69660
rect 7719 69600 7783 69604
rect 2584 69116 2648 69120
rect 2584 69060 2588 69116
rect 2588 69060 2644 69116
rect 2644 69060 2648 69116
rect 2584 69056 2648 69060
rect 2664 69116 2728 69120
rect 2664 69060 2668 69116
rect 2668 69060 2724 69116
rect 2724 69060 2728 69116
rect 2664 69056 2728 69060
rect 2744 69116 2808 69120
rect 2744 69060 2748 69116
rect 2748 69060 2804 69116
rect 2804 69060 2808 69116
rect 2744 69056 2808 69060
rect 2824 69116 2888 69120
rect 2824 69060 2828 69116
rect 2828 69060 2884 69116
rect 2884 69060 2888 69116
rect 2824 69056 2888 69060
rect 5847 69116 5911 69120
rect 5847 69060 5851 69116
rect 5851 69060 5907 69116
rect 5907 69060 5911 69116
rect 5847 69056 5911 69060
rect 5927 69116 5991 69120
rect 5927 69060 5931 69116
rect 5931 69060 5987 69116
rect 5987 69060 5991 69116
rect 5927 69056 5991 69060
rect 6007 69116 6071 69120
rect 6007 69060 6011 69116
rect 6011 69060 6067 69116
rect 6067 69060 6071 69116
rect 6007 69056 6071 69060
rect 6087 69116 6151 69120
rect 6087 69060 6091 69116
rect 6091 69060 6147 69116
rect 6147 69060 6151 69116
rect 6087 69056 6151 69060
rect 9111 69116 9175 69120
rect 9111 69060 9115 69116
rect 9115 69060 9171 69116
rect 9171 69060 9175 69116
rect 9111 69056 9175 69060
rect 9191 69116 9255 69120
rect 9191 69060 9195 69116
rect 9195 69060 9251 69116
rect 9251 69060 9255 69116
rect 9191 69056 9255 69060
rect 9271 69116 9335 69120
rect 9271 69060 9275 69116
rect 9275 69060 9331 69116
rect 9331 69060 9335 69116
rect 9271 69056 9335 69060
rect 9351 69116 9415 69120
rect 9351 69060 9355 69116
rect 9355 69060 9411 69116
rect 9411 69060 9415 69116
rect 9351 69056 9415 69060
rect 1716 68988 1780 69052
rect 2084 68580 2148 68644
rect 4215 68572 4279 68576
rect 4215 68516 4219 68572
rect 4219 68516 4275 68572
rect 4275 68516 4279 68572
rect 4215 68512 4279 68516
rect 4295 68572 4359 68576
rect 4295 68516 4299 68572
rect 4299 68516 4355 68572
rect 4355 68516 4359 68572
rect 4295 68512 4359 68516
rect 4375 68572 4439 68576
rect 4375 68516 4379 68572
rect 4379 68516 4435 68572
rect 4435 68516 4439 68572
rect 4375 68512 4439 68516
rect 4455 68572 4519 68576
rect 4455 68516 4459 68572
rect 4459 68516 4515 68572
rect 4515 68516 4519 68572
rect 4455 68512 4519 68516
rect 7479 68572 7543 68576
rect 7479 68516 7483 68572
rect 7483 68516 7539 68572
rect 7539 68516 7543 68572
rect 7479 68512 7543 68516
rect 7559 68572 7623 68576
rect 7559 68516 7563 68572
rect 7563 68516 7619 68572
rect 7619 68516 7623 68572
rect 7559 68512 7623 68516
rect 7639 68572 7703 68576
rect 7639 68516 7643 68572
rect 7643 68516 7699 68572
rect 7699 68516 7703 68572
rect 7639 68512 7703 68516
rect 7719 68572 7783 68576
rect 7719 68516 7723 68572
rect 7723 68516 7779 68572
rect 7779 68516 7783 68572
rect 7719 68512 7783 68516
rect 2584 68028 2648 68032
rect 2584 67972 2588 68028
rect 2588 67972 2644 68028
rect 2644 67972 2648 68028
rect 2584 67968 2648 67972
rect 2664 68028 2728 68032
rect 2664 67972 2668 68028
rect 2668 67972 2724 68028
rect 2724 67972 2728 68028
rect 2664 67968 2728 67972
rect 2744 68028 2808 68032
rect 2744 67972 2748 68028
rect 2748 67972 2804 68028
rect 2804 67972 2808 68028
rect 2744 67968 2808 67972
rect 2824 68028 2888 68032
rect 2824 67972 2828 68028
rect 2828 67972 2884 68028
rect 2884 67972 2888 68028
rect 2824 67968 2888 67972
rect 5847 68028 5911 68032
rect 5847 67972 5851 68028
rect 5851 67972 5907 68028
rect 5907 67972 5911 68028
rect 5847 67968 5911 67972
rect 5927 68028 5991 68032
rect 5927 67972 5931 68028
rect 5931 67972 5987 68028
rect 5987 67972 5991 68028
rect 5927 67968 5991 67972
rect 6007 68028 6071 68032
rect 6007 67972 6011 68028
rect 6011 67972 6067 68028
rect 6067 67972 6071 68028
rect 6007 67968 6071 67972
rect 6087 68028 6151 68032
rect 6087 67972 6091 68028
rect 6091 67972 6147 68028
rect 6147 67972 6151 68028
rect 6087 67968 6151 67972
rect 9111 68028 9175 68032
rect 9111 67972 9115 68028
rect 9115 67972 9171 68028
rect 9171 67972 9175 68028
rect 9111 67968 9175 67972
rect 9191 68028 9255 68032
rect 9191 67972 9195 68028
rect 9195 67972 9251 68028
rect 9251 67972 9255 68028
rect 9191 67968 9255 67972
rect 9271 68028 9335 68032
rect 9271 67972 9275 68028
rect 9275 67972 9331 68028
rect 9331 67972 9335 68028
rect 9271 67968 9335 67972
rect 9351 68028 9415 68032
rect 9351 67972 9355 68028
rect 9355 67972 9411 68028
rect 9411 67972 9415 68028
rect 9351 67968 9415 67972
rect 1532 67824 1596 67828
rect 1532 67768 1546 67824
rect 1546 67768 1596 67824
rect 1532 67764 1596 67768
rect 4215 67484 4279 67488
rect 4215 67428 4219 67484
rect 4219 67428 4275 67484
rect 4275 67428 4279 67484
rect 4215 67424 4279 67428
rect 4295 67484 4359 67488
rect 4295 67428 4299 67484
rect 4299 67428 4355 67484
rect 4355 67428 4359 67484
rect 4295 67424 4359 67428
rect 4375 67484 4439 67488
rect 4375 67428 4379 67484
rect 4379 67428 4435 67484
rect 4435 67428 4439 67484
rect 4375 67424 4439 67428
rect 4455 67484 4519 67488
rect 4455 67428 4459 67484
rect 4459 67428 4515 67484
rect 4515 67428 4519 67484
rect 4455 67424 4519 67428
rect 7479 67484 7543 67488
rect 7479 67428 7483 67484
rect 7483 67428 7539 67484
rect 7539 67428 7543 67484
rect 7479 67424 7543 67428
rect 7559 67484 7623 67488
rect 7559 67428 7563 67484
rect 7563 67428 7619 67484
rect 7619 67428 7623 67484
rect 7559 67424 7623 67428
rect 7639 67484 7703 67488
rect 7639 67428 7643 67484
rect 7643 67428 7699 67484
rect 7699 67428 7703 67484
rect 7639 67424 7703 67428
rect 7719 67484 7783 67488
rect 7719 67428 7723 67484
rect 7723 67428 7779 67484
rect 7779 67428 7783 67484
rect 7719 67424 7783 67428
rect 2584 66940 2648 66944
rect 2584 66884 2588 66940
rect 2588 66884 2644 66940
rect 2644 66884 2648 66940
rect 2584 66880 2648 66884
rect 2664 66940 2728 66944
rect 2664 66884 2668 66940
rect 2668 66884 2724 66940
rect 2724 66884 2728 66940
rect 2664 66880 2728 66884
rect 2744 66940 2808 66944
rect 2744 66884 2748 66940
rect 2748 66884 2804 66940
rect 2804 66884 2808 66940
rect 2744 66880 2808 66884
rect 2824 66940 2888 66944
rect 2824 66884 2828 66940
rect 2828 66884 2884 66940
rect 2884 66884 2888 66940
rect 2824 66880 2888 66884
rect 5847 66940 5911 66944
rect 5847 66884 5851 66940
rect 5851 66884 5907 66940
rect 5907 66884 5911 66940
rect 5847 66880 5911 66884
rect 5927 66940 5991 66944
rect 5927 66884 5931 66940
rect 5931 66884 5987 66940
rect 5987 66884 5991 66940
rect 5927 66880 5991 66884
rect 6007 66940 6071 66944
rect 6007 66884 6011 66940
rect 6011 66884 6067 66940
rect 6067 66884 6071 66940
rect 6007 66880 6071 66884
rect 6087 66940 6151 66944
rect 6087 66884 6091 66940
rect 6091 66884 6147 66940
rect 6147 66884 6151 66940
rect 6087 66880 6151 66884
rect 9111 66940 9175 66944
rect 9111 66884 9115 66940
rect 9115 66884 9171 66940
rect 9171 66884 9175 66940
rect 9111 66880 9175 66884
rect 9191 66940 9255 66944
rect 9191 66884 9195 66940
rect 9195 66884 9251 66940
rect 9251 66884 9255 66940
rect 9191 66880 9255 66884
rect 9271 66940 9335 66944
rect 9271 66884 9275 66940
rect 9275 66884 9331 66940
rect 9331 66884 9335 66940
rect 9271 66880 9335 66884
rect 9351 66940 9415 66944
rect 9351 66884 9355 66940
rect 9355 66884 9411 66940
rect 9411 66884 9415 66940
rect 9351 66880 9415 66884
rect 4215 66396 4279 66400
rect 4215 66340 4219 66396
rect 4219 66340 4275 66396
rect 4275 66340 4279 66396
rect 4215 66336 4279 66340
rect 4295 66396 4359 66400
rect 4295 66340 4299 66396
rect 4299 66340 4355 66396
rect 4355 66340 4359 66396
rect 4295 66336 4359 66340
rect 4375 66396 4439 66400
rect 4375 66340 4379 66396
rect 4379 66340 4435 66396
rect 4435 66340 4439 66396
rect 4375 66336 4439 66340
rect 4455 66396 4519 66400
rect 4455 66340 4459 66396
rect 4459 66340 4515 66396
rect 4515 66340 4519 66396
rect 4455 66336 4519 66340
rect 7479 66396 7543 66400
rect 7479 66340 7483 66396
rect 7483 66340 7539 66396
rect 7539 66340 7543 66396
rect 7479 66336 7543 66340
rect 7559 66396 7623 66400
rect 7559 66340 7563 66396
rect 7563 66340 7619 66396
rect 7619 66340 7623 66396
rect 7559 66336 7623 66340
rect 7639 66396 7703 66400
rect 7639 66340 7643 66396
rect 7643 66340 7699 66396
rect 7699 66340 7703 66396
rect 7639 66336 7703 66340
rect 7719 66396 7783 66400
rect 7719 66340 7723 66396
rect 7723 66340 7779 66396
rect 7779 66340 7783 66396
rect 7719 66336 7783 66340
rect 2584 65852 2648 65856
rect 2584 65796 2588 65852
rect 2588 65796 2644 65852
rect 2644 65796 2648 65852
rect 2584 65792 2648 65796
rect 2664 65852 2728 65856
rect 2664 65796 2668 65852
rect 2668 65796 2724 65852
rect 2724 65796 2728 65852
rect 2664 65792 2728 65796
rect 2744 65852 2808 65856
rect 2744 65796 2748 65852
rect 2748 65796 2804 65852
rect 2804 65796 2808 65852
rect 2744 65792 2808 65796
rect 2824 65852 2888 65856
rect 2824 65796 2828 65852
rect 2828 65796 2884 65852
rect 2884 65796 2888 65852
rect 2824 65792 2888 65796
rect 5847 65852 5911 65856
rect 5847 65796 5851 65852
rect 5851 65796 5907 65852
rect 5907 65796 5911 65852
rect 5847 65792 5911 65796
rect 5927 65852 5991 65856
rect 5927 65796 5931 65852
rect 5931 65796 5987 65852
rect 5987 65796 5991 65852
rect 5927 65792 5991 65796
rect 6007 65852 6071 65856
rect 6007 65796 6011 65852
rect 6011 65796 6067 65852
rect 6067 65796 6071 65852
rect 6007 65792 6071 65796
rect 6087 65852 6151 65856
rect 6087 65796 6091 65852
rect 6091 65796 6147 65852
rect 6147 65796 6151 65852
rect 6087 65792 6151 65796
rect 9111 65852 9175 65856
rect 9111 65796 9115 65852
rect 9115 65796 9171 65852
rect 9171 65796 9175 65852
rect 9111 65792 9175 65796
rect 9191 65852 9255 65856
rect 9191 65796 9195 65852
rect 9195 65796 9251 65852
rect 9251 65796 9255 65852
rect 9191 65792 9255 65796
rect 9271 65852 9335 65856
rect 9271 65796 9275 65852
rect 9275 65796 9331 65852
rect 9331 65796 9335 65852
rect 9271 65792 9335 65796
rect 9351 65852 9415 65856
rect 9351 65796 9355 65852
rect 9355 65796 9411 65852
rect 9411 65796 9415 65852
rect 9351 65792 9415 65796
rect 4215 65308 4279 65312
rect 4215 65252 4219 65308
rect 4219 65252 4275 65308
rect 4275 65252 4279 65308
rect 4215 65248 4279 65252
rect 4295 65308 4359 65312
rect 4295 65252 4299 65308
rect 4299 65252 4355 65308
rect 4355 65252 4359 65308
rect 4295 65248 4359 65252
rect 4375 65308 4439 65312
rect 4375 65252 4379 65308
rect 4379 65252 4435 65308
rect 4435 65252 4439 65308
rect 4375 65248 4439 65252
rect 4455 65308 4519 65312
rect 4455 65252 4459 65308
rect 4459 65252 4515 65308
rect 4515 65252 4519 65308
rect 4455 65248 4519 65252
rect 7479 65308 7543 65312
rect 7479 65252 7483 65308
rect 7483 65252 7539 65308
rect 7539 65252 7543 65308
rect 7479 65248 7543 65252
rect 7559 65308 7623 65312
rect 7559 65252 7563 65308
rect 7563 65252 7619 65308
rect 7619 65252 7623 65308
rect 7559 65248 7623 65252
rect 7639 65308 7703 65312
rect 7639 65252 7643 65308
rect 7643 65252 7699 65308
rect 7699 65252 7703 65308
rect 7639 65248 7703 65252
rect 7719 65308 7783 65312
rect 7719 65252 7723 65308
rect 7723 65252 7779 65308
rect 7779 65252 7783 65308
rect 7719 65248 7783 65252
rect 2268 64832 2332 64836
rect 2268 64776 2318 64832
rect 2318 64776 2332 64832
rect 2268 64772 2332 64776
rect 2584 64764 2648 64768
rect 2584 64708 2588 64764
rect 2588 64708 2644 64764
rect 2644 64708 2648 64764
rect 2584 64704 2648 64708
rect 2664 64764 2728 64768
rect 2664 64708 2668 64764
rect 2668 64708 2724 64764
rect 2724 64708 2728 64764
rect 2664 64704 2728 64708
rect 2744 64764 2808 64768
rect 2744 64708 2748 64764
rect 2748 64708 2804 64764
rect 2804 64708 2808 64764
rect 2744 64704 2808 64708
rect 2824 64764 2888 64768
rect 2824 64708 2828 64764
rect 2828 64708 2884 64764
rect 2884 64708 2888 64764
rect 2824 64704 2888 64708
rect 5847 64764 5911 64768
rect 5847 64708 5851 64764
rect 5851 64708 5907 64764
rect 5907 64708 5911 64764
rect 5847 64704 5911 64708
rect 5927 64764 5991 64768
rect 5927 64708 5931 64764
rect 5931 64708 5987 64764
rect 5987 64708 5991 64764
rect 5927 64704 5991 64708
rect 6007 64764 6071 64768
rect 6007 64708 6011 64764
rect 6011 64708 6067 64764
rect 6067 64708 6071 64764
rect 6007 64704 6071 64708
rect 6087 64764 6151 64768
rect 6087 64708 6091 64764
rect 6091 64708 6147 64764
rect 6147 64708 6151 64764
rect 6087 64704 6151 64708
rect 9111 64764 9175 64768
rect 9111 64708 9115 64764
rect 9115 64708 9171 64764
rect 9171 64708 9175 64764
rect 9111 64704 9175 64708
rect 9191 64764 9255 64768
rect 9191 64708 9195 64764
rect 9195 64708 9251 64764
rect 9251 64708 9255 64764
rect 9191 64704 9255 64708
rect 9271 64764 9335 64768
rect 9271 64708 9275 64764
rect 9275 64708 9331 64764
rect 9331 64708 9335 64764
rect 9271 64704 9335 64708
rect 9351 64764 9415 64768
rect 9351 64708 9355 64764
rect 9355 64708 9411 64764
rect 9411 64708 9415 64764
rect 9351 64704 9415 64708
rect 4215 64220 4279 64224
rect 4215 64164 4219 64220
rect 4219 64164 4275 64220
rect 4275 64164 4279 64220
rect 4215 64160 4279 64164
rect 4295 64220 4359 64224
rect 4295 64164 4299 64220
rect 4299 64164 4355 64220
rect 4355 64164 4359 64220
rect 4295 64160 4359 64164
rect 4375 64220 4439 64224
rect 4375 64164 4379 64220
rect 4379 64164 4435 64220
rect 4435 64164 4439 64220
rect 4375 64160 4439 64164
rect 4455 64220 4519 64224
rect 4455 64164 4459 64220
rect 4459 64164 4515 64220
rect 4515 64164 4519 64220
rect 4455 64160 4519 64164
rect 7479 64220 7543 64224
rect 7479 64164 7483 64220
rect 7483 64164 7539 64220
rect 7539 64164 7543 64220
rect 7479 64160 7543 64164
rect 7559 64220 7623 64224
rect 7559 64164 7563 64220
rect 7563 64164 7619 64220
rect 7619 64164 7623 64220
rect 7559 64160 7623 64164
rect 7639 64220 7703 64224
rect 7639 64164 7643 64220
rect 7643 64164 7699 64220
rect 7699 64164 7703 64220
rect 7639 64160 7703 64164
rect 7719 64220 7783 64224
rect 7719 64164 7723 64220
rect 7723 64164 7779 64220
rect 7779 64164 7783 64220
rect 7719 64160 7783 64164
rect 2584 63676 2648 63680
rect 2584 63620 2588 63676
rect 2588 63620 2644 63676
rect 2644 63620 2648 63676
rect 2584 63616 2648 63620
rect 2664 63676 2728 63680
rect 2664 63620 2668 63676
rect 2668 63620 2724 63676
rect 2724 63620 2728 63676
rect 2664 63616 2728 63620
rect 2744 63676 2808 63680
rect 2744 63620 2748 63676
rect 2748 63620 2804 63676
rect 2804 63620 2808 63676
rect 2744 63616 2808 63620
rect 2824 63676 2888 63680
rect 2824 63620 2828 63676
rect 2828 63620 2884 63676
rect 2884 63620 2888 63676
rect 2824 63616 2888 63620
rect 5847 63676 5911 63680
rect 5847 63620 5851 63676
rect 5851 63620 5907 63676
rect 5907 63620 5911 63676
rect 5847 63616 5911 63620
rect 5927 63676 5991 63680
rect 5927 63620 5931 63676
rect 5931 63620 5987 63676
rect 5987 63620 5991 63676
rect 5927 63616 5991 63620
rect 6007 63676 6071 63680
rect 6007 63620 6011 63676
rect 6011 63620 6067 63676
rect 6067 63620 6071 63676
rect 6007 63616 6071 63620
rect 6087 63676 6151 63680
rect 6087 63620 6091 63676
rect 6091 63620 6147 63676
rect 6147 63620 6151 63676
rect 6087 63616 6151 63620
rect 9111 63676 9175 63680
rect 9111 63620 9115 63676
rect 9115 63620 9171 63676
rect 9171 63620 9175 63676
rect 9111 63616 9175 63620
rect 9191 63676 9255 63680
rect 9191 63620 9195 63676
rect 9195 63620 9251 63676
rect 9251 63620 9255 63676
rect 9191 63616 9255 63620
rect 9271 63676 9335 63680
rect 9271 63620 9275 63676
rect 9275 63620 9331 63676
rect 9331 63620 9335 63676
rect 9271 63616 9335 63620
rect 9351 63676 9415 63680
rect 9351 63620 9355 63676
rect 9355 63620 9411 63676
rect 9411 63620 9415 63676
rect 9351 63616 9415 63620
rect 4215 63132 4279 63136
rect 4215 63076 4219 63132
rect 4219 63076 4275 63132
rect 4275 63076 4279 63132
rect 4215 63072 4279 63076
rect 4295 63132 4359 63136
rect 4295 63076 4299 63132
rect 4299 63076 4355 63132
rect 4355 63076 4359 63132
rect 4295 63072 4359 63076
rect 4375 63132 4439 63136
rect 4375 63076 4379 63132
rect 4379 63076 4435 63132
rect 4435 63076 4439 63132
rect 4375 63072 4439 63076
rect 4455 63132 4519 63136
rect 4455 63076 4459 63132
rect 4459 63076 4515 63132
rect 4515 63076 4519 63132
rect 4455 63072 4519 63076
rect 7479 63132 7543 63136
rect 7479 63076 7483 63132
rect 7483 63076 7539 63132
rect 7539 63076 7543 63132
rect 7479 63072 7543 63076
rect 7559 63132 7623 63136
rect 7559 63076 7563 63132
rect 7563 63076 7619 63132
rect 7619 63076 7623 63132
rect 7559 63072 7623 63076
rect 7639 63132 7703 63136
rect 7639 63076 7643 63132
rect 7643 63076 7699 63132
rect 7699 63076 7703 63132
rect 7639 63072 7703 63076
rect 7719 63132 7783 63136
rect 7719 63076 7723 63132
rect 7723 63076 7779 63132
rect 7779 63076 7783 63132
rect 7719 63072 7783 63076
rect 2584 62588 2648 62592
rect 2584 62532 2588 62588
rect 2588 62532 2644 62588
rect 2644 62532 2648 62588
rect 2584 62528 2648 62532
rect 2664 62588 2728 62592
rect 2664 62532 2668 62588
rect 2668 62532 2724 62588
rect 2724 62532 2728 62588
rect 2664 62528 2728 62532
rect 2744 62588 2808 62592
rect 2744 62532 2748 62588
rect 2748 62532 2804 62588
rect 2804 62532 2808 62588
rect 2744 62528 2808 62532
rect 2824 62588 2888 62592
rect 2824 62532 2828 62588
rect 2828 62532 2884 62588
rect 2884 62532 2888 62588
rect 2824 62528 2888 62532
rect 5847 62588 5911 62592
rect 5847 62532 5851 62588
rect 5851 62532 5907 62588
rect 5907 62532 5911 62588
rect 5847 62528 5911 62532
rect 5927 62588 5991 62592
rect 5927 62532 5931 62588
rect 5931 62532 5987 62588
rect 5987 62532 5991 62588
rect 5927 62528 5991 62532
rect 6007 62588 6071 62592
rect 6007 62532 6011 62588
rect 6011 62532 6067 62588
rect 6067 62532 6071 62588
rect 6007 62528 6071 62532
rect 6087 62588 6151 62592
rect 6087 62532 6091 62588
rect 6091 62532 6147 62588
rect 6147 62532 6151 62588
rect 6087 62528 6151 62532
rect 9111 62588 9175 62592
rect 9111 62532 9115 62588
rect 9115 62532 9171 62588
rect 9171 62532 9175 62588
rect 9111 62528 9175 62532
rect 9191 62588 9255 62592
rect 9191 62532 9195 62588
rect 9195 62532 9251 62588
rect 9251 62532 9255 62588
rect 9191 62528 9255 62532
rect 9271 62588 9335 62592
rect 9271 62532 9275 62588
rect 9275 62532 9331 62588
rect 9331 62532 9335 62588
rect 9271 62528 9335 62532
rect 9351 62588 9415 62592
rect 9351 62532 9355 62588
rect 9355 62532 9411 62588
rect 9411 62532 9415 62588
rect 9351 62528 9415 62532
rect 2084 62052 2148 62116
rect 4215 62044 4279 62048
rect 4215 61988 4219 62044
rect 4219 61988 4275 62044
rect 4275 61988 4279 62044
rect 4215 61984 4279 61988
rect 4295 62044 4359 62048
rect 4295 61988 4299 62044
rect 4299 61988 4355 62044
rect 4355 61988 4359 62044
rect 4295 61984 4359 61988
rect 4375 62044 4439 62048
rect 4375 61988 4379 62044
rect 4379 61988 4435 62044
rect 4435 61988 4439 62044
rect 4375 61984 4439 61988
rect 4455 62044 4519 62048
rect 4455 61988 4459 62044
rect 4459 61988 4515 62044
rect 4515 61988 4519 62044
rect 4455 61984 4519 61988
rect 7479 62044 7543 62048
rect 7479 61988 7483 62044
rect 7483 61988 7539 62044
rect 7539 61988 7543 62044
rect 7479 61984 7543 61988
rect 7559 62044 7623 62048
rect 7559 61988 7563 62044
rect 7563 61988 7619 62044
rect 7619 61988 7623 62044
rect 7559 61984 7623 61988
rect 7639 62044 7703 62048
rect 7639 61988 7643 62044
rect 7643 61988 7699 62044
rect 7699 61988 7703 62044
rect 7639 61984 7703 61988
rect 7719 62044 7783 62048
rect 7719 61988 7723 62044
rect 7723 61988 7779 62044
rect 7779 61988 7783 62044
rect 7719 61984 7783 61988
rect 2268 61508 2332 61572
rect 2584 61500 2648 61504
rect 2584 61444 2588 61500
rect 2588 61444 2644 61500
rect 2644 61444 2648 61500
rect 2584 61440 2648 61444
rect 2664 61500 2728 61504
rect 2664 61444 2668 61500
rect 2668 61444 2724 61500
rect 2724 61444 2728 61500
rect 2664 61440 2728 61444
rect 2744 61500 2808 61504
rect 2744 61444 2748 61500
rect 2748 61444 2804 61500
rect 2804 61444 2808 61500
rect 2744 61440 2808 61444
rect 2824 61500 2888 61504
rect 2824 61444 2828 61500
rect 2828 61444 2884 61500
rect 2884 61444 2888 61500
rect 2824 61440 2888 61444
rect 5847 61500 5911 61504
rect 5847 61444 5851 61500
rect 5851 61444 5907 61500
rect 5907 61444 5911 61500
rect 5847 61440 5911 61444
rect 5927 61500 5991 61504
rect 5927 61444 5931 61500
rect 5931 61444 5987 61500
rect 5987 61444 5991 61500
rect 5927 61440 5991 61444
rect 6007 61500 6071 61504
rect 6007 61444 6011 61500
rect 6011 61444 6067 61500
rect 6067 61444 6071 61500
rect 6007 61440 6071 61444
rect 6087 61500 6151 61504
rect 6087 61444 6091 61500
rect 6091 61444 6147 61500
rect 6147 61444 6151 61500
rect 6087 61440 6151 61444
rect 9111 61500 9175 61504
rect 9111 61444 9115 61500
rect 9115 61444 9171 61500
rect 9171 61444 9175 61500
rect 9111 61440 9175 61444
rect 9191 61500 9255 61504
rect 9191 61444 9195 61500
rect 9195 61444 9251 61500
rect 9251 61444 9255 61500
rect 9191 61440 9255 61444
rect 9271 61500 9335 61504
rect 9271 61444 9275 61500
rect 9275 61444 9331 61500
rect 9331 61444 9335 61500
rect 9271 61440 9335 61444
rect 9351 61500 9415 61504
rect 9351 61444 9355 61500
rect 9355 61444 9411 61500
rect 9411 61444 9415 61500
rect 9351 61440 9415 61444
rect 4215 60956 4279 60960
rect 4215 60900 4219 60956
rect 4219 60900 4275 60956
rect 4275 60900 4279 60956
rect 4215 60896 4279 60900
rect 4295 60956 4359 60960
rect 4295 60900 4299 60956
rect 4299 60900 4355 60956
rect 4355 60900 4359 60956
rect 4295 60896 4359 60900
rect 4375 60956 4439 60960
rect 4375 60900 4379 60956
rect 4379 60900 4435 60956
rect 4435 60900 4439 60956
rect 4375 60896 4439 60900
rect 4455 60956 4519 60960
rect 4455 60900 4459 60956
rect 4459 60900 4515 60956
rect 4515 60900 4519 60956
rect 4455 60896 4519 60900
rect 7479 60956 7543 60960
rect 7479 60900 7483 60956
rect 7483 60900 7539 60956
rect 7539 60900 7543 60956
rect 7479 60896 7543 60900
rect 7559 60956 7623 60960
rect 7559 60900 7563 60956
rect 7563 60900 7619 60956
rect 7619 60900 7623 60956
rect 7559 60896 7623 60900
rect 7639 60956 7703 60960
rect 7639 60900 7643 60956
rect 7643 60900 7699 60956
rect 7699 60900 7703 60956
rect 7639 60896 7703 60900
rect 7719 60956 7783 60960
rect 7719 60900 7723 60956
rect 7723 60900 7779 60956
rect 7779 60900 7783 60956
rect 7719 60896 7783 60900
rect 2584 60412 2648 60416
rect 2584 60356 2588 60412
rect 2588 60356 2644 60412
rect 2644 60356 2648 60412
rect 2584 60352 2648 60356
rect 2664 60412 2728 60416
rect 2664 60356 2668 60412
rect 2668 60356 2724 60412
rect 2724 60356 2728 60412
rect 2664 60352 2728 60356
rect 2744 60412 2808 60416
rect 2744 60356 2748 60412
rect 2748 60356 2804 60412
rect 2804 60356 2808 60412
rect 2744 60352 2808 60356
rect 2824 60412 2888 60416
rect 2824 60356 2828 60412
rect 2828 60356 2884 60412
rect 2884 60356 2888 60412
rect 2824 60352 2888 60356
rect 5847 60412 5911 60416
rect 5847 60356 5851 60412
rect 5851 60356 5907 60412
rect 5907 60356 5911 60412
rect 5847 60352 5911 60356
rect 5927 60412 5991 60416
rect 5927 60356 5931 60412
rect 5931 60356 5987 60412
rect 5987 60356 5991 60412
rect 5927 60352 5991 60356
rect 6007 60412 6071 60416
rect 6007 60356 6011 60412
rect 6011 60356 6067 60412
rect 6067 60356 6071 60412
rect 6007 60352 6071 60356
rect 6087 60412 6151 60416
rect 6087 60356 6091 60412
rect 6091 60356 6147 60412
rect 6147 60356 6151 60412
rect 6087 60352 6151 60356
rect 9111 60412 9175 60416
rect 9111 60356 9115 60412
rect 9115 60356 9171 60412
rect 9171 60356 9175 60412
rect 9111 60352 9175 60356
rect 9191 60412 9255 60416
rect 9191 60356 9195 60412
rect 9195 60356 9251 60412
rect 9251 60356 9255 60412
rect 9191 60352 9255 60356
rect 9271 60412 9335 60416
rect 9271 60356 9275 60412
rect 9275 60356 9331 60412
rect 9331 60356 9335 60412
rect 9271 60352 9335 60356
rect 9351 60412 9415 60416
rect 9351 60356 9355 60412
rect 9355 60356 9411 60412
rect 9411 60356 9415 60412
rect 9351 60352 9415 60356
rect 4215 59868 4279 59872
rect 4215 59812 4219 59868
rect 4219 59812 4275 59868
rect 4275 59812 4279 59868
rect 4215 59808 4279 59812
rect 4295 59868 4359 59872
rect 4295 59812 4299 59868
rect 4299 59812 4355 59868
rect 4355 59812 4359 59868
rect 4295 59808 4359 59812
rect 4375 59868 4439 59872
rect 4375 59812 4379 59868
rect 4379 59812 4435 59868
rect 4435 59812 4439 59868
rect 4375 59808 4439 59812
rect 4455 59868 4519 59872
rect 4455 59812 4459 59868
rect 4459 59812 4515 59868
rect 4515 59812 4519 59868
rect 4455 59808 4519 59812
rect 7479 59868 7543 59872
rect 7479 59812 7483 59868
rect 7483 59812 7539 59868
rect 7539 59812 7543 59868
rect 7479 59808 7543 59812
rect 7559 59868 7623 59872
rect 7559 59812 7563 59868
rect 7563 59812 7619 59868
rect 7619 59812 7623 59868
rect 7559 59808 7623 59812
rect 7639 59868 7703 59872
rect 7639 59812 7643 59868
rect 7643 59812 7699 59868
rect 7699 59812 7703 59868
rect 7639 59808 7703 59812
rect 7719 59868 7783 59872
rect 7719 59812 7723 59868
rect 7723 59812 7779 59868
rect 7779 59812 7783 59868
rect 7719 59808 7783 59812
rect 2584 59324 2648 59328
rect 2584 59268 2588 59324
rect 2588 59268 2644 59324
rect 2644 59268 2648 59324
rect 2584 59264 2648 59268
rect 2664 59324 2728 59328
rect 2664 59268 2668 59324
rect 2668 59268 2724 59324
rect 2724 59268 2728 59324
rect 2664 59264 2728 59268
rect 2744 59324 2808 59328
rect 2744 59268 2748 59324
rect 2748 59268 2804 59324
rect 2804 59268 2808 59324
rect 2744 59264 2808 59268
rect 2824 59324 2888 59328
rect 2824 59268 2828 59324
rect 2828 59268 2884 59324
rect 2884 59268 2888 59324
rect 2824 59264 2888 59268
rect 5847 59324 5911 59328
rect 5847 59268 5851 59324
rect 5851 59268 5907 59324
rect 5907 59268 5911 59324
rect 5847 59264 5911 59268
rect 5927 59324 5991 59328
rect 5927 59268 5931 59324
rect 5931 59268 5987 59324
rect 5987 59268 5991 59324
rect 5927 59264 5991 59268
rect 6007 59324 6071 59328
rect 6007 59268 6011 59324
rect 6011 59268 6067 59324
rect 6067 59268 6071 59324
rect 6007 59264 6071 59268
rect 6087 59324 6151 59328
rect 6087 59268 6091 59324
rect 6091 59268 6147 59324
rect 6147 59268 6151 59324
rect 6087 59264 6151 59268
rect 9111 59324 9175 59328
rect 9111 59268 9115 59324
rect 9115 59268 9171 59324
rect 9171 59268 9175 59324
rect 9111 59264 9175 59268
rect 9191 59324 9255 59328
rect 9191 59268 9195 59324
rect 9195 59268 9251 59324
rect 9251 59268 9255 59324
rect 9191 59264 9255 59268
rect 9271 59324 9335 59328
rect 9271 59268 9275 59324
rect 9275 59268 9331 59324
rect 9331 59268 9335 59324
rect 9271 59264 9335 59268
rect 9351 59324 9415 59328
rect 9351 59268 9355 59324
rect 9355 59268 9411 59324
rect 9411 59268 9415 59324
rect 9351 59264 9415 59268
rect 4215 58780 4279 58784
rect 4215 58724 4219 58780
rect 4219 58724 4275 58780
rect 4275 58724 4279 58780
rect 4215 58720 4279 58724
rect 4295 58780 4359 58784
rect 4295 58724 4299 58780
rect 4299 58724 4355 58780
rect 4355 58724 4359 58780
rect 4295 58720 4359 58724
rect 4375 58780 4439 58784
rect 4375 58724 4379 58780
rect 4379 58724 4435 58780
rect 4435 58724 4439 58780
rect 4375 58720 4439 58724
rect 4455 58780 4519 58784
rect 4455 58724 4459 58780
rect 4459 58724 4515 58780
rect 4515 58724 4519 58780
rect 4455 58720 4519 58724
rect 7479 58780 7543 58784
rect 7479 58724 7483 58780
rect 7483 58724 7539 58780
rect 7539 58724 7543 58780
rect 7479 58720 7543 58724
rect 7559 58780 7623 58784
rect 7559 58724 7563 58780
rect 7563 58724 7619 58780
rect 7619 58724 7623 58780
rect 7559 58720 7623 58724
rect 7639 58780 7703 58784
rect 7639 58724 7643 58780
rect 7643 58724 7699 58780
rect 7699 58724 7703 58780
rect 7639 58720 7703 58724
rect 7719 58780 7783 58784
rect 7719 58724 7723 58780
rect 7723 58724 7779 58780
rect 7779 58724 7783 58780
rect 7719 58720 7783 58724
rect 1716 58304 1780 58308
rect 1716 58248 1730 58304
rect 1730 58248 1780 58304
rect 1716 58244 1780 58248
rect 2584 58236 2648 58240
rect 2584 58180 2588 58236
rect 2588 58180 2644 58236
rect 2644 58180 2648 58236
rect 2584 58176 2648 58180
rect 2664 58236 2728 58240
rect 2664 58180 2668 58236
rect 2668 58180 2724 58236
rect 2724 58180 2728 58236
rect 2664 58176 2728 58180
rect 2744 58236 2808 58240
rect 2744 58180 2748 58236
rect 2748 58180 2804 58236
rect 2804 58180 2808 58236
rect 2744 58176 2808 58180
rect 2824 58236 2888 58240
rect 2824 58180 2828 58236
rect 2828 58180 2884 58236
rect 2884 58180 2888 58236
rect 2824 58176 2888 58180
rect 5847 58236 5911 58240
rect 5847 58180 5851 58236
rect 5851 58180 5907 58236
rect 5907 58180 5911 58236
rect 5847 58176 5911 58180
rect 5927 58236 5991 58240
rect 5927 58180 5931 58236
rect 5931 58180 5987 58236
rect 5987 58180 5991 58236
rect 5927 58176 5991 58180
rect 6007 58236 6071 58240
rect 6007 58180 6011 58236
rect 6011 58180 6067 58236
rect 6067 58180 6071 58236
rect 6007 58176 6071 58180
rect 6087 58236 6151 58240
rect 6087 58180 6091 58236
rect 6091 58180 6147 58236
rect 6147 58180 6151 58236
rect 6087 58176 6151 58180
rect 9111 58236 9175 58240
rect 9111 58180 9115 58236
rect 9115 58180 9171 58236
rect 9171 58180 9175 58236
rect 9111 58176 9175 58180
rect 9191 58236 9255 58240
rect 9191 58180 9195 58236
rect 9195 58180 9251 58236
rect 9251 58180 9255 58236
rect 9191 58176 9255 58180
rect 9271 58236 9335 58240
rect 9271 58180 9275 58236
rect 9275 58180 9331 58236
rect 9331 58180 9335 58236
rect 9271 58176 9335 58180
rect 9351 58236 9415 58240
rect 9351 58180 9355 58236
rect 9355 58180 9411 58236
rect 9411 58180 9415 58236
rect 9351 58176 9415 58180
rect 4215 57692 4279 57696
rect 4215 57636 4219 57692
rect 4219 57636 4275 57692
rect 4275 57636 4279 57692
rect 4215 57632 4279 57636
rect 4295 57692 4359 57696
rect 4295 57636 4299 57692
rect 4299 57636 4355 57692
rect 4355 57636 4359 57692
rect 4295 57632 4359 57636
rect 4375 57692 4439 57696
rect 4375 57636 4379 57692
rect 4379 57636 4435 57692
rect 4435 57636 4439 57692
rect 4375 57632 4439 57636
rect 4455 57692 4519 57696
rect 4455 57636 4459 57692
rect 4459 57636 4515 57692
rect 4515 57636 4519 57692
rect 4455 57632 4519 57636
rect 7479 57692 7543 57696
rect 7479 57636 7483 57692
rect 7483 57636 7539 57692
rect 7539 57636 7543 57692
rect 7479 57632 7543 57636
rect 7559 57692 7623 57696
rect 7559 57636 7563 57692
rect 7563 57636 7619 57692
rect 7619 57636 7623 57692
rect 7559 57632 7623 57636
rect 7639 57692 7703 57696
rect 7639 57636 7643 57692
rect 7643 57636 7699 57692
rect 7699 57636 7703 57692
rect 7639 57632 7703 57636
rect 7719 57692 7783 57696
rect 7719 57636 7723 57692
rect 7723 57636 7779 57692
rect 7779 57636 7783 57692
rect 7719 57632 7783 57636
rect 2584 57148 2648 57152
rect 2584 57092 2588 57148
rect 2588 57092 2644 57148
rect 2644 57092 2648 57148
rect 2584 57088 2648 57092
rect 2664 57148 2728 57152
rect 2664 57092 2668 57148
rect 2668 57092 2724 57148
rect 2724 57092 2728 57148
rect 2664 57088 2728 57092
rect 2744 57148 2808 57152
rect 2744 57092 2748 57148
rect 2748 57092 2804 57148
rect 2804 57092 2808 57148
rect 2744 57088 2808 57092
rect 2824 57148 2888 57152
rect 2824 57092 2828 57148
rect 2828 57092 2884 57148
rect 2884 57092 2888 57148
rect 2824 57088 2888 57092
rect 5847 57148 5911 57152
rect 5847 57092 5851 57148
rect 5851 57092 5907 57148
rect 5907 57092 5911 57148
rect 5847 57088 5911 57092
rect 5927 57148 5991 57152
rect 5927 57092 5931 57148
rect 5931 57092 5987 57148
rect 5987 57092 5991 57148
rect 5927 57088 5991 57092
rect 6007 57148 6071 57152
rect 6007 57092 6011 57148
rect 6011 57092 6067 57148
rect 6067 57092 6071 57148
rect 6007 57088 6071 57092
rect 6087 57148 6151 57152
rect 6087 57092 6091 57148
rect 6091 57092 6147 57148
rect 6147 57092 6151 57148
rect 6087 57088 6151 57092
rect 9111 57148 9175 57152
rect 9111 57092 9115 57148
rect 9115 57092 9171 57148
rect 9171 57092 9175 57148
rect 9111 57088 9175 57092
rect 9191 57148 9255 57152
rect 9191 57092 9195 57148
rect 9195 57092 9251 57148
rect 9251 57092 9255 57148
rect 9191 57088 9255 57092
rect 9271 57148 9335 57152
rect 9271 57092 9275 57148
rect 9275 57092 9331 57148
rect 9331 57092 9335 57148
rect 9271 57088 9335 57092
rect 9351 57148 9415 57152
rect 9351 57092 9355 57148
rect 9355 57092 9411 57148
rect 9411 57092 9415 57148
rect 9351 57088 9415 57092
rect 3004 56672 3068 56676
rect 3004 56616 3054 56672
rect 3054 56616 3068 56672
rect 3004 56612 3068 56616
rect 4215 56604 4279 56608
rect 4215 56548 4219 56604
rect 4219 56548 4275 56604
rect 4275 56548 4279 56604
rect 4215 56544 4279 56548
rect 4295 56604 4359 56608
rect 4295 56548 4299 56604
rect 4299 56548 4355 56604
rect 4355 56548 4359 56604
rect 4295 56544 4359 56548
rect 4375 56604 4439 56608
rect 4375 56548 4379 56604
rect 4379 56548 4435 56604
rect 4435 56548 4439 56604
rect 4375 56544 4439 56548
rect 4455 56604 4519 56608
rect 4455 56548 4459 56604
rect 4459 56548 4515 56604
rect 4515 56548 4519 56604
rect 4455 56544 4519 56548
rect 7479 56604 7543 56608
rect 7479 56548 7483 56604
rect 7483 56548 7539 56604
rect 7539 56548 7543 56604
rect 7479 56544 7543 56548
rect 7559 56604 7623 56608
rect 7559 56548 7563 56604
rect 7563 56548 7619 56604
rect 7619 56548 7623 56604
rect 7559 56544 7623 56548
rect 7639 56604 7703 56608
rect 7639 56548 7643 56604
rect 7643 56548 7699 56604
rect 7699 56548 7703 56604
rect 7639 56544 7703 56548
rect 7719 56604 7783 56608
rect 7719 56548 7723 56604
rect 7723 56548 7779 56604
rect 7779 56548 7783 56604
rect 7719 56544 7783 56548
rect 4660 56204 4724 56268
rect 2584 56060 2648 56064
rect 2584 56004 2588 56060
rect 2588 56004 2644 56060
rect 2644 56004 2648 56060
rect 2584 56000 2648 56004
rect 2664 56060 2728 56064
rect 2664 56004 2668 56060
rect 2668 56004 2724 56060
rect 2724 56004 2728 56060
rect 2664 56000 2728 56004
rect 2744 56060 2808 56064
rect 2744 56004 2748 56060
rect 2748 56004 2804 56060
rect 2804 56004 2808 56060
rect 2744 56000 2808 56004
rect 2824 56060 2888 56064
rect 2824 56004 2828 56060
rect 2828 56004 2884 56060
rect 2884 56004 2888 56060
rect 2824 56000 2888 56004
rect 5847 56060 5911 56064
rect 5847 56004 5851 56060
rect 5851 56004 5907 56060
rect 5907 56004 5911 56060
rect 5847 56000 5911 56004
rect 5927 56060 5991 56064
rect 5927 56004 5931 56060
rect 5931 56004 5987 56060
rect 5987 56004 5991 56060
rect 5927 56000 5991 56004
rect 6007 56060 6071 56064
rect 6007 56004 6011 56060
rect 6011 56004 6067 56060
rect 6067 56004 6071 56060
rect 6007 56000 6071 56004
rect 6087 56060 6151 56064
rect 6087 56004 6091 56060
rect 6091 56004 6147 56060
rect 6147 56004 6151 56060
rect 6087 56000 6151 56004
rect 9111 56060 9175 56064
rect 9111 56004 9115 56060
rect 9115 56004 9171 56060
rect 9171 56004 9175 56060
rect 9111 56000 9175 56004
rect 9191 56060 9255 56064
rect 9191 56004 9195 56060
rect 9195 56004 9251 56060
rect 9251 56004 9255 56060
rect 9191 56000 9255 56004
rect 9271 56060 9335 56064
rect 9271 56004 9275 56060
rect 9275 56004 9331 56060
rect 9331 56004 9335 56060
rect 9271 56000 9335 56004
rect 9351 56060 9415 56064
rect 9351 56004 9355 56060
rect 9355 56004 9411 56060
rect 9411 56004 9415 56060
rect 9351 56000 9415 56004
rect 3188 55796 3252 55860
rect 4215 55516 4279 55520
rect 4215 55460 4219 55516
rect 4219 55460 4275 55516
rect 4275 55460 4279 55516
rect 4215 55456 4279 55460
rect 4295 55516 4359 55520
rect 4295 55460 4299 55516
rect 4299 55460 4355 55516
rect 4355 55460 4359 55516
rect 4295 55456 4359 55460
rect 4375 55516 4439 55520
rect 4375 55460 4379 55516
rect 4379 55460 4435 55516
rect 4435 55460 4439 55516
rect 4375 55456 4439 55460
rect 4455 55516 4519 55520
rect 4455 55460 4459 55516
rect 4459 55460 4515 55516
rect 4515 55460 4519 55516
rect 4455 55456 4519 55460
rect 7479 55516 7543 55520
rect 7479 55460 7483 55516
rect 7483 55460 7539 55516
rect 7539 55460 7543 55516
rect 7479 55456 7543 55460
rect 7559 55516 7623 55520
rect 7559 55460 7563 55516
rect 7563 55460 7619 55516
rect 7619 55460 7623 55516
rect 7559 55456 7623 55460
rect 7639 55516 7703 55520
rect 7639 55460 7643 55516
rect 7643 55460 7699 55516
rect 7699 55460 7703 55516
rect 7639 55456 7703 55460
rect 7719 55516 7783 55520
rect 7719 55460 7723 55516
rect 7723 55460 7779 55516
rect 7779 55460 7783 55516
rect 7719 55456 7783 55460
rect 1164 55252 1228 55316
rect 2584 54972 2648 54976
rect 2584 54916 2588 54972
rect 2588 54916 2644 54972
rect 2644 54916 2648 54972
rect 2584 54912 2648 54916
rect 2664 54972 2728 54976
rect 2664 54916 2668 54972
rect 2668 54916 2724 54972
rect 2724 54916 2728 54972
rect 2664 54912 2728 54916
rect 2744 54972 2808 54976
rect 2744 54916 2748 54972
rect 2748 54916 2804 54972
rect 2804 54916 2808 54972
rect 2744 54912 2808 54916
rect 2824 54972 2888 54976
rect 2824 54916 2828 54972
rect 2828 54916 2884 54972
rect 2884 54916 2888 54972
rect 2824 54912 2888 54916
rect 5847 54972 5911 54976
rect 5847 54916 5851 54972
rect 5851 54916 5907 54972
rect 5907 54916 5911 54972
rect 5847 54912 5911 54916
rect 5927 54972 5991 54976
rect 5927 54916 5931 54972
rect 5931 54916 5987 54972
rect 5987 54916 5991 54972
rect 5927 54912 5991 54916
rect 6007 54972 6071 54976
rect 6007 54916 6011 54972
rect 6011 54916 6067 54972
rect 6067 54916 6071 54972
rect 6007 54912 6071 54916
rect 6087 54972 6151 54976
rect 6087 54916 6091 54972
rect 6091 54916 6147 54972
rect 6147 54916 6151 54972
rect 6087 54912 6151 54916
rect 9111 54972 9175 54976
rect 9111 54916 9115 54972
rect 9115 54916 9171 54972
rect 9171 54916 9175 54972
rect 9111 54912 9175 54916
rect 9191 54972 9255 54976
rect 9191 54916 9195 54972
rect 9195 54916 9251 54972
rect 9251 54916 9255 54972
rect 9191 54912 9255 54916
rect 9271 54972 9335 54976
rect 9271 54916 9275 54972
rect 9275 54916 9331 54972
rect 9331 54916 9335 54972
rect 9271 54912 9335 54916
rect 9351 54972 9415 54976
rect 9351 54916 9355 54972
rect 9355 54916 9411 54972
rect 9411 54916 9415 54972
rect 9351 54912 9415 54916
rect 3372 54708 3436 54772
rect 4215 54428 4279 54432
rect 4215 54372 4219 54428
rect 4219 54372 4275 54428
rect 4275 54372 4279 54428
rect 4215 54368 4279 54372
rect 4295 54428 4359 54432
rect 4295 54372 4299 54428
rect 4299 54372 4355 54428
rect 4355 54372 4359 54428
rect 4295 54368 4359 54372
rect 4375 54428 4439 54432
rect 4375 54372 4379 54428
rect 4379 54372 4435 54428
rect 4435 54372 4439 54428
rect 4375 54368 4439 54372
rect 4455 54428 4519 54432
rect 4455 54372 4459 54428
rect 4459 54372 4515 54428
rect 4515 54372 4519 54428
rect 4455 54368 4519 54372
rect 7479 54428 7543 54432
rect 7479 54372 7483 54428
rect 7483 54372 7539 54428
rect 7539 54372 7543 54428
rect 7479 54368 7543 54372
rect 7559 54428 7623 54432
rect 7559 54372 7563 54428
rect 7563 54372 7619 54428
rect 7619 54372 7623 54428
rect 7559 54368 7623 54372
rect 7639 54428 7703 54432
rect 7639 54372 7643 54428
rect 7643 54372 7699 54428
rect 7699 54372 7703 54428
rect 7639 54368 7703 54372
rect 7719 54428 7783 54432
rect 7719 54372 7723 54428
rect 7723 54372 7779 54428
rect 7779 54372 7783 54428
rect 7719 54368 7783 54372
rect 2584 53884 2648 53888
rect 2584 53828 2588 53884
rect 2588 53828 2644 53884
rect 2644 53828 2648 53884
rect 2584 53824 2648 53828
rect 2664 53884 2728 53888
rect 2664 53828 2668 53884
rect 2668 53828 2724 53884
rect 2724 53828 2728 53884
rect 2664 53824 2728 53828
rect 2744 53884 2808 53888
rect 2744 53828 2748 53884
rect 2748 53828 2804 53884
rect 2804 53828 2808 53884
rect 2744 53824 2808 53828
rect 2824 53884 2888 53888
rect 2824 53828 2828 53884
rect 2828 53828 2884 53884
rect 2884 53828 2888 53884
rect 2824 53824 2888 53828
rect 5847 53884 5911 53888
rect 5847 53828 5851 53884
rect 5851 53828 5907 53884
rect 5907 53828 5911 53884
rect 5847 53824 5911 53828
rect 5927 53884 5991 53888
rect 5927 53828 5931 53884
rect 5931 53828 5987 53884
rect 5987 53828 5991 53884
rect 5927 53824 5991 53828
rect 6007 53884 6071 53888
rect 6007 53828 6011 53884
rect 6011 53828 6067 53884
rect 6067 53828 6071 53884
rect 6007 53824 6071 53828
rect 6087 53884 6151 53888
rect 6087 53828 6091 53884
rect 6091 53828 6147 53884
rect 6147 53828 6151 53884
rect 6087 53824 6151 53828
rect 9111 53884 9175 53888
rect 9111 53828 9115 53884
rect 9115 53828 9171 53884
rect 9171 53828 9175 53884
rect 9111 53824 9175 53828
rect 9191 53884 9255 53888
rect 9191 53828 9195 53884
rect 9195 53828 9251 53884
rect 9251 53828 9255 53884
rect 9191 53824 9255 53828
rect 9271 53884 9335 53888
rect 9271 53828 9275 53884
rect 9275 53828 9331 53884
rect 9331 53828 9335 53884
rect 9271 53824 9335 53828
rect 9351 53884 9415 53888
rect 9351 53828 9355 53884
rect 9355 53828 9411 53884
rect 9411 53828 9415 53884
rect 9351 53824 9415 53828
rect 5396 53680 5460 53684
rect 5396 53624 5446 53680
rect 5446 53624 5460 53680
rect 5396 53620 5460 53624
rect 2268 53348 2332 53412
rect 4215 53340 4279 53344
rect 4215 53284 4219 53340
rect 4219 53284 4275 53340
rect 4275 53284 4279 53340
rect 4215 53280 4279 53284
rect 4295 53340 4359 53344
rect 4295 53284 4299 53340
rect 4299 53284 4355 53340
rect 4355 53284 4359 53340
rect 4295 53280 4359 53284
rect 4375 53340 4439 53344
rect 4375 53284 4379 53340
rect 4379 53284 4435 53340
rect 4435 53284 4439 53340
rect 4375 53280 4439 53284
rect 4455 53340 4519 53344
rect 4455 53284 4459 53340
rect 4459 53284 4515 53340
rect 4515 53284 4519 53340
rect 4455 53280 4519 53284
rect 7479 53340 7543 53344
rect 7479 53284 7483 53340
rect 7483 53284 7539 53340
rect 7539 53284 7543 53340
rect 7479 53280 7543 53284
rect 7559 53340 7623 53344
rect 7559 53284 7563 53340
rect 7563 53284 7619 53340
rect 7619 53284 7623 53340
rect 7559 53280 7623 53284
rect 7639 53340 7703 53344
rect 7639 53284 7643 53340
rect 7643 53284 7699 53340
rect 7699 53284 7703 53340
rect 7639 53280 7703 53284
rect 7719 53340 7783 53344
rect 7719 53284 7723 53340
rect 7723 53284 7779 53340
rect 7779 53284 7783 53340
rect 7719 53280 7783 53284
rect 4844 53076 4908 53140
rect 2584 52796 2648 52800
rect 2584 52740 2588 52796
rect 2588 52740 2644 52796
rect 2644 52740 2648 52796
rect 2584 52736 2648 52740
rect 2664 52796 2728 52800
rect 2664 52740 2668 52796
rect 2668 52740 2724 52796
rect 2724 52740 2728 52796
rect 2664 52736 2728 52740
rect 2744 52796 2808 52800
rect 2744 52740 2748 52796
rect 2748 52740 2804 52796
rect 2804 52740 2808 52796
rect 2744 52736 2808 52740
rect 2824 52796 2888 52800
rect 2824 52740 2828 52796
rect 2828 52740 2884 52796
rect 2884 52740 2888 52796
rect 2824 52736 2888 52740
rect 5847 52796 5911 52800
rect 5847 52740 5851 52796
rect 5851 52740 5907 52796
rect 5907 52740 5911 52796
rect 5847 52736 5911 52740
rect 5927 52796 5991 52800
rect 5927 52740 5931 52796
rect 5931 52740 5987 52796
rect 5987 52740 5991 52796
rect 5927 52736 5991 52740
rect 6007 52796 6071 52800
rect 6007 52740 6011 52796
rect 6011 52740 6067 52796
rect 6067 52740 6071 52796
rect 6007 52736 6071 52740
rect 6087 52796 6151 52800
rect 6087 52740 6091 52796
rect 6091 52740 6147 52796
rect 6147 52740 6151 52796
rect 6087 52736 6151 52740
rect 9111 52796 9175 52800
rect 9111 52740 9115 52796
rect 9115 52740 9171 52796
rect 9171 52740 9175 52796
rect 9111 52736 9175 52740
rect 9191 52796 9255 52800
rect 9191 52740 9195 52796
rect 9195 52740 9251 52796
rect 9251 52740 9255 52796
rect 9191 52736 9255 52740
rect 9271 52796 9335 52800
rect 9271 52740 9275 52796
rect 9275 52740 9331 52796
rect 9331 52740 9335 52796
rect 9271 52736 9335 52740
rect 9351 52796 9415 52800
rect 9351 52740 9355 52796
rect 9355 52740 9411 52796
rect 9411 52740 9415 52796
rect 9351 52736 9415 52740
rect 4215 52252 4279 52256
rect 4215 52196 4219 52252
rect 4219 52196 4275 52252
rect 4275 52196 4279 52252
rect 4215 52192 4279 52196
rect 4295 52252 4359 52256
rect 4295 52196 4299 52252
rect 4299 52196 4355 52252
rect 4355 52196 4359 52252
rect 4295 52192 4359 52196
rect 4375 52252 4439 52256
rect 4375 52196 4379 52252
rect 4379 52196 4435 52252
rect 4435 52196 4439 52252
rect 4375 52192 4439 52196
rect 4455 52252 4519 52256
rect 4455 52196 4459 52252
rect 4459 52196 4515 52252
rect 4515 52196 4519 52252
rect 4455 52192 4519 52196
rect 7479 52252 7543 52256
rect 7479 52196 7483 52252
rect 7483 52196 7539 52252
rect 7539 52196 7543 52252
rect 7479 52192 7543 52196
rect 7559 52252 7623 52256
rect 7559 52196 7563 52252
rect 7563 52196 7619 52252
rect 7619 52196 7623 52252
rect 7559 52192 7623 52196
rect 7639 52252 7703 52256
rect 7639 52196 7643 52252
rect 7643 52196 7699 52252
rect 7699 52196 7703 52252
rect 7639 52192 7703 52196
rect 7719 52252 7783 52256
rect 7719 52196 7723 52252
rect 7723 52196 7779 52252
rect 7779 52196 7783 52252
rect 7719 52192 7783 52196
rect 2584 51708 2648 51712
rect 2584 51652 2588 51708
rect 2588 51652 2644 51708
rect 2644 51652 2648 51708
rect 2584 51648 2648 51652
rect 2664 51708 2728 51712
rect 2664 51652 2668 51708
rect 2668 51652 2724 51708
rect 2724 51652 2728 51708
rect 2664 51648 2728 51652
rect 2744 51708 2808 51712
rect 2744 51652 2748 51708
rect 2748 51652 2804 51708
rect 2804 51652 2808 51708
rect 2744 51648 2808 51652
rect 2824 51708 2888 51712
rect 2824 51652 2828 51708
rect 2828 51652 2884 51708
rect 2884 51652 2888 51708
rect 2824 51648 2888 51652
rect 5847 51708 5911 51712
rect 5847 51652 5851 51708
rect 5851 51652 5907 51708
rect 5907 51652 5911 51708
rect 5847 51648 5911 51652
rect 5927 51708 5991 51712
rect 5927 51652 5931 51708
rect 5931 51652 5987 51708
rect 5987 51652 5991 51708
rect 5927 51648 5991 51652
rect 6007 51708 6071 51712
rect 6007 51652 6011 51708
rect 6011 51652 6067 51708
rect 6067 51652 6071 51708
rect 6007 51648 6071 51652
rect 6087 51708 6151 51712
rect 6087 51652 6091 51708
rect 6091 51652 6147 51708
rect 6147 51652 6151 51708
rect 6087 51648 6151 51652
rect 9111 51708 9175 51712
rect 9111 51652 9115 51708
rect 9115 51652 9171 51708
rect 9171 51652 9175 51708
rect 9111 51648 9175 51652
rect 9191 51708 9255 51712
rect 9191 51652 9195 51708
rect 9195 51652 9251 51708
rect 9251 51652 9255 51708
rect 9191 51648 9255 51652
rect 9271 51708 9335 51712
rect 9271 51652 9275 51708
rect 9275 51652 9331 51708
rect 9331 51652 9335 51708
rect 9271 51648 9335 51652
rect 9351 51708 9415 51712
rect 9351 51652 9355 51708
rect 9355 51652 9411 51708
rect 9411 51652 9415 51708
rect 9351 51648 9415 51652
rect 4844 51640 4908 51644
rect 4844 51584 4858 51640
rect 4858 51584 4908 51640
rect 4844 51580 4908 51584
rect 2268 51232 2332 51236
rect 2268 51176 2318 51232
rect 2318 51176 2332 51232
rect 2268 51172 2332 51176
rect 4215 51164 4279 51168
rect 4215 51108 4219 51164
rect 4219 51108 4275 51164
rect 4275 51108 4279 51164
rect 4215 51104 4279 51108
rect 4295 51164 4359 51168
rect 4295 51108 4299 51164
rect 4299 51108 4355 51164
rect 4355 51108 4359 51164
rect 4295 51104 4359 51108
rect 4375 51164 4439 51168
rect 4375 51108 4379 51164
rect 4379 51108 4435 51164
rect 4435 51108 4439 51164
rect 4375 51104 4439 51108
rect 4455 51164 4519 51168
rect 4455 51108 4459 51164
rect 4459 51108 4515 51164
rect 4515 51108 4519 51164
rect 4455 51104 4519 51108
rect 7479 51164 7543 51168
rect 7479 51108 7483 51164
rect 7483 51108 7539 51164
rect 7539 51108 7543 51164
rect 7479 51104 7543 51108
rect 7559 51164 7623 51168
rect 7559 51108 7563 51164
rect 7563 51108 7619 51164
rect 7619 51108 7623 51164
rect 7559 51104 7623 51108
rect 7639 51164 7703 51168
rect 7639 51108 7643 51164
rect 7643 51108 7699 51164
rect 7699 51108 7703 51164
rect 7639 51104 7703 51108
rect 7719 51164 7783 51168
rect 7719 51108 7723 51164
rect 7723 51108 7779 51164
rect 7779 51108 7783 51164
rect 7719 51104 7783 51108
rect 5396 51096 5460 51100
rect 5396 51040 5446 51096
rect 5446 51040 5460 51096
rect 5396 51036 5460 51040
rect 3188 50628 3252 50692
rect 2584 50620 2648 50624
rect 2584 50564 2588 50620
rect 2588 50564 2644 50620
rect 2644 50564 2648 50620
rect 2584 50560 2648 50564
rect 2664 50620 2728 50624
rect 2664 50564 2668 50620
rect 2668 50564 2724 50620
rect 2724 50564 2728 50620
rect 2664 50560 2728 50564
rect 2744 50620 2808 50624
rect 2744 50564 2748 50620
rect 2748 50564 2804 50620
rect 2804 50564 2808 50620
rect 2744 50560 2808 50564
rect 2824 50620 2888 50624
rect 2824 50564 2828 50620
rect 2828 50564 2884 50620
rect 2884 50564 2888 50620
rect 2824 50560 2888 50564
rect 5847 50620 5911 50624
rect 5847 50564 5851 50620
rect 5851 50564 5907 50620
rect 5907 50564 5911 50620
rect 5847 50560 5911 50564
rect 5927 50620 5991 50624
rect 5927 50564 5931 50620
rect 5931 50564 5987 50620
rect 5987 50564 5991 50620
rect 5927 50560 5991 50564
rect 6007 50620 6071 50624
rect 6007 50564 6011 50620
rect 6011 50564 6067 50620
rect 6067 50564 6071 50620
rect 6007 50560 6071 50564
rect 6087 50620 6151 50624
rect 6087 50564 6091 50620
rect 6091 50564 6147 50620
rect 6147 50564 6151 50620
rect 6087 50560 6151 50564
rect 9111 50620 9175 50624
rect 9111 50564 9115 50620
rect 9115 50564 9171 50620
rect 9171 50564 9175 50620
rect 9111 50560 9175 50564
rect 9191 50620 9255 50624
rect 9191 50564 9195 50620
rect 9195 50564 9251 50620
rect 9251 50564 9255 50620
rect 9191 50560 9255 50564
rect 9271 50620 9335 50624
rect 9271 50564 9275 50620
rect 9275 50564 9331 50620
rect 9331 50564 9335 50620
rect 9271 50560 9335 50564
rect 9351 50620 9415 50624
rect 9351 50564 9355 50620
rect 9355 50564 9411 50620
rect 9411 50564 9415 50620
rect 9351 50560 9415 50564
rect 4215 50076 4279 50080
rect 4215 50020 4219 50076
rect 4219 50020 4275 50076
rect 4275 50020 4279 50076
rect 4215 50016 4279 50020
rect 4295 50076 4359 50080
rect 4295 50020 4299 50076
rect 4299 50020 4355 50076
rect 4355 50020 4359 50076
rect 4295 50016 4359 50020
rect 4375 50076 4439 50080
rect 4375 50020 4379 50076
rect 4379 50020 4435 50076
rect 4435 50020 4439 50076
rect 4375 50016 4439 50020
rect 4455 50076 4519 50080
rect 4455 50020 4459 50076
rect 4459 50020 4515 50076
rect 4515 50020 4519 50076
rect 4455 50016 4519 50020
rect 7479 50076 7543 50080
rect 7479 50020 7483 50076
rect 7483 50020 7539 50076
rect 7539 50020 7543 50076
rect 7479 50016 7543 50020
rect 7559 50076 7623 50080
rect 7559 50020 7563 50076
rect 7563 50020 7619 50076
rect 7619 50020 7623 50076
rect 7559 50016 7623 50020
rect 7639 50076 7703 50080
rect 7639 50020 7643 50076
rect 7643 50020 7699 50076
rect 7699 50020 7703 50076
rect 7639 50016 7703 50020
rect 7719 50076 7783 50080
rect 7719 50020 7723 50076
rect 7723 50020 7779 50076
rect 7779 50020 7783 50076
rect 7719 50016 7783 50020
rect 2584 49532 2648 49536
rect 2584 49476 2588 49532
rect 2588 49476 2644 49532
rect 2644 49476 2648 49532
rect 2584 49472 2648 49476
rect 2664 49532 2728 49536
rect 2664 49476 2668 49532
rect 2668 49476 2724 49532
rect 2724 49476 2728 49532
rect 2664 49472 2728 49476
rect 2744 49532 2808 49536
rect 2744 49476 2748 49532
rect 2748 49476 2804 49532
rect 2804 49476 2808 49532
rect 2744 49472 2808 49476
rect 2824 49532 2888 49536
rect 2824 49476 2828 49532
rect 2828 49476 2884 49532
rect 2884 49476 2888 49532
rect 2824 49472 2888 49476
rect 5847 49532 5911 49536
rect 5847 49476 5851 49532
rect 5851 49476 5907 49532
rect 5907 49476 5911 49532
rect 5847 49472 5911 49476
rect 5927 49532 5991 49536
rect 5927 49476 5931 49532
rect 5931 49476 5987 49532
rect 5987 49476 5991 49532
rect 5927 49472 5991 49476
rect 6007 49532 6071 49536
rect 6007 49476 6011 49532
rect 6011 49476 6067 49532
rect 6067 49476 6071 49532
rect 6007 49472 6071 49476
rect 6087 49532 6151 49536
rect 6087 49476 6091 49532
rect 6091 49476 6147 49532
rect 6147 49476 6151 49532
rect 6087 49472 6151 49476
rect 9111 49532 9175 49536
rect 9111 49476 9115 49532
rect 9115 49476 9171 49532
rect 9171 49476 9175 49532
rect 9111 49472 9175 49476
rect 9191 49532 9255 49536
rect 9191 49476 9195 49532
rect 9195 49476 9251 49532
rect 9251 49476 9255 49532
rect 9191 49472 9255 49476
rect 9271 49532 9335 49536
rect 9271 49476 9275 49532
rect 9275 49476 9331 49532
rect 9331 49476 9335 49532
rect 9271 49472 9335 49476
rect 9351 49532 9415 49536
rect 9351 49476 9355 49532
rect 9355 49476 9411 49532
rect 9411 49476 9415 49532
rect 9351 49472 9415 49476
rect 3372 49268 3436 49332
rect 4215 48988 4279 48992
rect 4215 48932 4219 48988
rect 4219 48932 4275 48988
rect 4275 48932 4279 48988
rect 4215 48928 4279 48932
rect 4295 48988 4359 48992
rect 4295 48932 4299 48988
rect 4299 48932 4355 48988
rect 4355 48932 4359 48988
rect 4295 48928 4359 48932
rect 4375 48988 4439 48992
rect 4375 48932 4379 48988
rect 4379 48932 4435 48988
rect 4435 48932 4439 48988
rect 4375 48928 4439 48932
rect 4455 48988 4519 48992
rect 4455 48932 4459 48988
rect 4459 48932 4515 48988
rect 4515 48932 4519 48988
rect 4455 48928 4519 48932
rect 7479 48988 7543 48992
rect 7479 48932 7483 48988
rect 7483 48932 7539 48988
rect 7539 48932 7543 48988
rect 7479 48928 7543 48932
rect 7559 48988 7623 48992
rect 7559 48932 7563 48988
rect 7563 48932 7619 48988
rect 7619 48932 7623 48988
rect 7559 48928 7623 48932
rect 7639 48988 7703 48992
rect 7639 48932 7643 48988
rect 7643 48932 7699 48988
rect 7699 48932 7703 48988
rect 7639 48928 7703 48932
rect 7719 48988 7783 48992
rect 7719 48932 7723 48988
rect 7723 48932 7779 48988
rect 7779 48932 7783 48988
rect 7719 48928 7783 48932
rect 4660 48724 4724 48788
rect 6684 48724 6748 48788
rect 2584 48444 2648 48448
rect 2584 48388 2588 48444
rect 2588 48388 2644 48444
rect 2644 48388 2648 48444
rect 2584 48384 2648 48388
rect 2664 48444 2728 48448
rect 2664 48388 2668 48444
rect 2668 48388 2724 48444
rect 2724 48388 2728 48444
rect 2664 48384 2728 48388
rect 2744 48444 2808 48448
rect 2744 48388 2748 48444
rect 2748 48388 2804 48444
rect 2804 48388 2808 48444
rect 2744 48384 2808 48388
rect 2824 48444 2888 48448
rect 2824 48388 2828 48444
rect 2828 48388 2884 48444
rect 2884 48388 2888 48444
rect 2824 48384 2888 48388
rect 5847 48444 5911 48448
rect 5847 48388 5851 48444
rect 5851 48388 5907 48444
rect 5907 48388 5911 48444
rect 5847 48384 5911 48388
rect 5927 48444 5991 48448
rect 5927 48388 5931 48444
rect 5931 48388 5987 48444
rect 5987 48388 5991 48444
rect 5927 48384 5991 48388
rect 6007 48444 6071 48448
rect 6007 48388 6011 48444
rect 6011 48388 6067 48444
rect 6067 48388 6071 48444
rect 6007 48384 6071 48388
rect 6087 48444 6151 48448
rect 6087 48388 6091 48444
rect 6091 48388 6147 48444
rect 6147 48388 6151 48444
rect 6087 48384 6151 48388
rect 9111 48444 9175 48448
rect 9111 48388 9115 48444
rect 9115 48388 9171 48444
rect 9171 48388 9175 48444
rect 9111 48384 9175 48388
rect 9191 48444 9255 48448
rect 9191 48388 9195 48444
rect 9195 48388 9251 48444
rect 9251 48388 9255 48444
rect 9191 48384 9255 48388
rect 9271 48444 9335 48448
rect 9271 48388 9275 48444
rect 9275 48388 9331 48444
rect 9331 48388 9335 48444
rect 9271 48384 9335 48388
rect 9351 48444 9415 48448
rect 9351 48388 9355 48444
rect 9355 48388 9411 48444
rect 9411 48388 9415 48444
rect 9351 48384 9415 48388
rect 3740 48180 3804 48244
rect 4660 48044 4724 48108
rect 4215 47900 4279 47904
rect 4215 47844 4219 47900
rect 4219 47844 4275 47900
rect 4275 47844 4279 47900
rect 4215 47840 4279 47844
rect 4295 47900 4359 47904
rect 4295 47844 4299 47900
rect 4299 47844 4355 47900
rect 4355 47844 4359 47900
rect 4295 47840 4359 47844
rect 4375 47900 4439 47904
rect 4375 47844 4379 47900
rect 4379 47844 4435 47900
rect 4435 47844 4439 47900
rect 4375 47840 4439 47844
rect 4455 47900 4519 47904
rect 4455 47844 4459 47900
rect 4459 47844 4515 47900
rect 4515 47844 4519 47900
rect 4455 47840 4519 47844
rect 7479 47900 7543 47904
rect 7479 47844 7483 47900
rect 7483 47844 7539 47900
rect 7539 47844 7543 47900
rect 7479 47840 7543 47844
rect 7559 47900 7623 47904
rect 7559 47844 7563 47900
rect 7563 47844 7619 47900
rect 7619 47844 7623 47900
rect 7559 47840 7623 47844
rect 7639 47900 7703 47904
rect 7639 47844 7643 47900
rect 7643 47844 7699 47900
rect 7699 47844 7703 47900
rect 7639 47840 7703 47844
rect 7719 47900 7783 47904
rect 7719 47844 7723 47900
rect 7723 47844 7779 47900
rect 7779 47844 7783 47900
rect 7719 47840 7783 47844
rect 2584 47356 2648 47360
rect 2584 47300 2588 47356
rect 2588 47300 2644 47356
rect 2644 47300 2648 47356
rect 2584 47296 2648 47300
rect 2664 47356 2728 47360
rect 2664 47300 2668 47356
rect 2668 47300 2724 47356
rect 2724 47300 2728 47356
rect 2664 47296 2728 47300
rect 2744 47356 2808 47360
rect 2744 47300 2748 47356
rect 2748 47300 2804 47356
rect 2804 47300 2808 47356
rect 2744 47296 2808 47300
rect 2824 47356 2888 47360
rect 2824 47300 2828 47356
rect 2828 47300 2884 47356
rect 2884 47300 2888 47356
rect 2824 47296 2888 47300
rect 5847 47356 5911 47360
rect 5847 47300 5851 47356
rect 5851 47300 5907 47356
rect 5907 47300 5911 47356
rect 5847 47296 5911 47300
rect 5927 47356 5991 47360
rect 5927 47300 5931 47356
rect 5931 47300 5987 47356
rect 5987 47300 5991 47356
rect 5927 47296 5991 47300
rect 6007 47356 6071 47360
rect 6007 47300 6011 47356
rect 6011 47300 6067 47356
rect 6067 47300 6071 47356
rect 6007 47296 6071 47300
rect 6087 47356 6151 47360
rect 6087 47300 6091 47356
rect 6091 47300 6147 47356
rect 6147 47300 6151 47356
rect 6087 47296 6151 47300
rect 9111 47356 9175 47360
rect 9111 47300 9115 47356
rect 9115 47300 9171 47356
rect 9171 47300 9175 47356
rect 9111 47296 9175 47300
rect 9191 47356 9255 47360
rect 9191 47300 9195 47356
rect 9195 47300 9251 47356
rect 9251 47300 9255 47356
rect 9191 47296 9255 47300
rect 9271 47356 9335 47360
rect 9271 47300 9275 47356
rect 9275 47300 9331 47356
rect 9331 47300 9335 47356
rect 9271 47296 9335 47300
rect 9351 47356 9415 47360
rect 9351 47300 9355 47356
rect 9355 47300 9411 47356
rect 9411 47300 9415 47356
rect 9351 47296 9415 47300
rect 3004 46820 3068 46884
rect 4215 46812 4279 46816
rect 4215 46756 4219 46812
rect 4219 46756 4275 46812
rect 4275 46756 4279 46812
rect 4215 46752 4279 46756
rect 4295 46812 4359 46816
rect 4295 46756 4299 46812
rect 4299 46756 4355 46812
rect 4355 46756 4359 46812
rect 4295 46752 4359 46756
rect 4375 46812 4439 46816
rect 4375 46756 4379 46812
rect 4379 46756 4435 46812
rect 4435 46756 4439 46812
rect 4375 46752 4439 46756
rect 4455 46812 4519 46816
rect 4455 46756 4459 46812
rect 4459 46756 4515 46812
rect 4515 46756 4519 46812
rect 4455 46752 4519 46756
rect 7479 46812 7543 46816
rect 7479 46756 7483 46812
rect 7483 46756 7539 46812
rect 7539 46756 7543 46812
rect 7479 46752 7543 46756
rect 7559 46812 7623 46816
rect 7559 46756 7563 46812
rect 7563 46756 7619 46812
rect 7619 46756 7623 46812
rect 7559 46752 7623 46756
rect 7639 46812 7703 46816
rect 7639 46756 7643 46812
rect 7643 46756 7699 46812
rect 7699 46756 7703 46812
rect 7639 46752 7703 46756
rect 7719 46812 7783 46816
rect 7719 46756 7723 46812
rect 7723 46756 7779 46812
rect 7779 46756 7783 46812
rect 7719 46752 7783 46756
rect 6684 46336 6748 46340
rect 6684 46280 6734 46336
rect 6734 46280 6748 46336
rect 6684 46276 6748 46280
rect 2584 46268 2648 46272
rect 2584 46212 2588 46268
rect 2588 46212 2644 46268
rect 2644 46212 2648 46268
rect 2584 46208 2648 46212
rect 2664 46268 2728 46272
rect 2664 46212 2668 46268
rect 2668 46212 2724 46268
rect 2724 46212 2728 46268
rect 2664 46208 2728 46212
rect 2744 46268 2808 46272
rect 2744 46212 2748 46268
rect 2748 46212 2804 46268
rect 2804 46212 2808 46268
rect 2744 46208 2808 46212
rect 2824 46268 2888 46272
rect 2824 46212 2828 46268
rect 2828 46212 2884 46268
rect 2884 46212 2888 46268
rect 2824 46208 2888 46212
rect 5847 46268 5911 46272
rect 5847 46212 5851 46268
rect 5851 46212 5907 46268
rect 5907 46212 5911 46268
rect 5847 46208 5911 46212
rect 5927 46268 5991 46272
rect 5927 46212 5931 46268
rect 5931 46212 5987 46268
rect 5987 46212 5991 46268
rect 5927 46208 5991 46212
rect 6007 46268 6071 46272
rect 6007 46212 6011 46268
rect 6011 46212 6067 46268
rect 6067 46212 6071 46268
rect 6007 46208 6071 46212
rect 6087 46268 6151 46272
rect 6087 46212 6091 46268
rect 6091 46212 6147 46268
rect 6147 46212 6151 46268
rect 6087 46208 6151 46212
rect 9111 46268 9175 46272
rect 9111 46212 9115 46268
rect 9115 46212 9171 46268
rect 9171 46212 9175 46268
rect 9111 46208 9175 46212
rect 9191 46268 9255 46272
rect 9191 46212 9195 46268
rect 9195 46212 9251 46268
rect 9251 46212 9255 46268
rect 9191 46208 9255 46212
rect 9271 46268 9335 46272
rect 9271 46212 9275 46268
rect 9275 46212 9331 46268
rect 9331 46212 9335 46268
rect 9271 46208 9335 46212
rect 9351 46268 9415 46272
rect 9351 46212 9355 46268
rect 9355 46212 9411 46268
rect 9411 46212 9415 46268
rect 9351 46208 9415 46212
rect 2268 46004 2332 46068
rect 4215 45724 4279 45728
rect 4215 45668 4219 45724
rect 4219 45668 4275 45724
rect 4275 45668 4279 45724
rect 4215 45664 4279 45668
rect 4295 45724 4359 45728
rect 4295 45668 4299 45724
rect 4299 45668 4355 45724
rect 4355 45668 4359 45724
rect 4295 45664 4359 45668
rect 4375 45724 4439 45728
rect 4375 45668 4379 45724
rect 4379 45668 4435 45724
rect 4435 45668 4439 45724
rect 4375 45664 4439 45668
rect 4455 45724 4519 45728
rect 4455 45668 4459 45724
rect 4459 45668 4515 45724
rect 4515 45668 4519 45724
rect 4455 45664 4519 45668
rect 7479 45724 7543 45728
rect 7479 45668 7483 45724
rect 7483 45668 7539 45724
rect 7539 45668 7543 45724
rect 7479 45664 7543 45668
rect 7559 45724 7623 45728
rect 7559 45668 7563 45724
rect 7563 45668 7619 45724
rect 7619 45668 7623 45724
rect 7559 45664 7623 45668
rect 7639 45724 7703 45728
rect 7639 45668 7643 45724
rect 7643 45668 7699 45724
rect 7699 45668 7703 45724
rect 7639 45664 7703 45668
rect 7719 45724 7783 45728
rect 7719 45668 7723 45724
rect 7723 45668 7779 45724
rect 7779 45668 7783 45724
rect 7719 45664 7783 45668
rect 2584 45180 2648 45184
rect 2584 45124 2588 45180
rect 2588 45124 2644 45180
rect 2644 45124 2648 45180
rect 2584 45120 2648 45124
rect 2664 45180 2728 45184
rect 2664 45124 2668 45180
rect 2668 45124 2724 45180
rect 2724 45124 2728 45180
rect 2664 45120 2728 45124
rect 2744 45180 2808 45184
rect 2744 45124 2748 45180
rect 2748 45124 2804 45180
rect 2804 45124 2808 45180
rect 2744 45120 2808 45124
rect 2824 45180 2888 45184
rect 2824 45124 2828 45180
rect 2828 45124 2884 45180
rect 2884 45124 2888 45180
rect 2824 45120 2888 45124
rect 5847 45180 5911 45184
rect 5847 45124 5851 45180
rect 5851 45124 5907 45180
rect 5907 45124 5911 45180
rect 5847 45120 5911 45124
rect 5927 45180 5991 45184
rect 5927 45124 5931 45180
rect 5931 45124 5987 45180
rect 5987 45124 5991 45180
rect 5927 45120 5991 45124
rect 6007 45180 6071 45184
rect 6007 45124 6011 45180
rect 6011 45124 6067 45180
rect 6067 45124 6071 45180
rect 6007 45120 6071 45124
rect 6087 45180 6151 45184
rect 6087 45124 6091 45180
rect 6091 45124 6147 45180
rect 6147 45124 6151 45180
rect 6087 45120 6151 45124
rect 9111 45180 9175 45184
rect 9111 45124 9115 45180
rect 9115 45124 9171 45180
rect 9171 45124 9175 45180
rect 9111 45120 9175 45124
rect 9191 45180 9255 45184
rect 9191 45124 9195 45180
rect 9195 45124 9251 45180
rect 9251 45124 9255 45180
rect 9191 45120 9255 45124
rect 9271 45180 9335 45184
rect 9271 45124 9275 45180
rect 9275 45124 9331 45180
rect 9331 45124 9335 45180
rect 9271 45120 9335 45124
rect 9351 45180 9415 45184
rect 9351 45124 9355 45180
rect 9355 45124 9411 45180
rect 9411 45124 9415 45180
rect 9351 45120 9415 45124
rect 4215 44636 4279 44640
rect 4215 44580 4219 44636
rect 4219 44580 4275 44636
rect 4275 44580 4279 44636
rect 4215 44576 4279 44580
rect 4295 44636 4359 44640
rect 4295 44580 4299 44636
rect 4299 44580 4355 44636
rect 4355 44580 4359 44636
rect 4295 44576 4359 44580
rect 4375 44636 4439 44640
rect 4375 44580 4379 44636
rect 4379 44580 4435 44636
rect 4435 44580 4439 44636
rect 4375 44576 4439 44580
rect 4455 44636 4519 44640
rect 4455 44580 4459 44636
rect 4459 44580 4515 44636
rect 4515 44580 4519 44636
rect 4455 44576 4519 44580
rect 7479 44636 7543 44640
rect 7479 44580 7483 44636
rect 7483 44580 7539 44636
rect 7539 44580 7543 44636
rect 7479 44576 7543 44580
rect 7559 44636 7623 44640
rect 7559 44580 7563 44636
rect 7563 44580 7619 44636
rect 7619 44580 7623 44636
rect 7559 44576 7623 44580
rect 7639 44636 7703 44640
rect 7639 44580 7643 44636
rect 7643 44580 7699 44636
rect 7699 44580 7703 44636
rect 7639 44576 7703 44580
rect 7719 44636 7783 44640
rect 7719 44580 7723 44636
rect 7723 44580 7779 44636
rect 7779 44580 7783 44636
rect 7719 44576 7783 44580
rect 2584 44092 2648 44096
rect 2584 44036 2588 44092
rect 2588 44036 2644 44092
rect 2644 44036 2648 44092
rect 2584 44032 2648 44036
rect 2664 44092 2728 44096
rect 2664 44036 2668 44092
rect 2668 44036 2724 44092
rect 2724 44036 2728 44092
rect 2664 44032 2728 44036
rect 2744 44092 2808 44096
rect 2744 44036 2748 44092
rect 2748 44036 2804 44092
rect 2804 44036 2808 44092
rect 2744 44032 2808 44036
rect 2824 44092 2888 44096
rect 2824 44036 2828 44092
rect 2828 44036 2884 44092
rect 2884 44036 2888 44092
rect 2824 44032 2888 44036
rect 5847 44092 5911 44096
rect 5847 44036 5851 44092
rect 5851 44036 5907 44092
rect 5907 44036 5911 44092
rect 5847 44032 5911 44036
rect 5927 44092 5991 44096
rect 5927 44036 5931 44092
rect 5931 44036 5987 44092
rect 5987 44036 5991 44092
rect 5927 44032 5991 44036
rect 6007 44092 6071 44096
rect 6007 44036 6011 44092
rect 6011 44036 6067 44092
rect 6067 44036 6071 44092
rect 6007 44032 6071 44036
rect 6087 44092 6151 44096
rect 6087 44036 6091 44092
rect 6091 44036 6147 44092
rect 6147 44036 6151 44092
rect 6087 44032 6151 44036
rect 9111 44092 9175 44096
rect 9111 44036 9115 44092
rect 9115 44036 9171 44092
rect 9171 44036 9175 44092
rect 9111 44032 9175 44036
rect 9191 44092 9255 44096
rect 9191 44036 9195 44092
rect 9195 44036 9251 44092
rect 9251 44036 9255 44092
rect 9191 44032 9255 44036
rect 9271 44092 9335 44096
rect 9271 44036 9275 44092
rect 9275 44036 9331 44092
rect 9331 44036 9335 44092
rect 9271 44032 9335 44036
rect 9351 44092 9415 44096
rect 9351 44036 9355 44092
rect 9355 44036 9411 44092
rect 9411 44036 9415 44092
rect 9351 44032 9415 44036
rect 4215 43548 4279 43552
rect 4215 43492 4219 43548
rect 4219 43492 4275 43548
rect 4275 43492 4279 43548
rect 4215 43488 4279 43492
rect 4295 43548 4359 43552
rect 4295 43492 4299 43548
rect 4299 43492 4355 43548
rect 4355 43492 4359 43548
rect 4295 43488 4359 43492
rect 4375 43548 4439 43552
rect 4375 43492 4379 43548
rect 4379 43492 4435 43548
rect 4435 43492 4439 43548
rect 4375 43488 4439 43492
rect 4455 43548 4519 43552
rect 4455 43492 4459 43548
rect 4459 43492 4515 43548
rect 4515 43492 4519 43548
rect 4455 43488 4519 43492
rect 7479 43548 7543 43552
rect 7479 43492 7483 43548
rect 7483 43492 7539 43548
rect 7539 43492 7543 43548
rect 7479 43488 7543 43492
rect 7559 43548 7623 43552
rect 7559 43492 7563 43548
rect 7563 43492 7619 43548
rect 7619 43492 7623 43548
rect 7559 43488 7623 43492
rect 7639 43548 7703 43552
rect 7639 43492 7643 43548
rect 7643 43492 7699 43548
rect 7699 43492 7703 43548
rect 7639 43488 7703 43492
rect 7719 43548 7783 43552
rect 7719 43492 7723 43548
rect 7723 43492 7779 43548
rect 7779 43492 7783 43548
rect 7719 43488 7783 43492
rect 3740 43148 3804 43212
rect 2584 43004 2648 43008
rect 2584 42948 2588 43004
rect 2588 42948 2644 43004
rect 2644 42948 2648 43004
rect 2584 42944 2648 42948
rect 2664 43004 2728 43008
rect 2664 42948 2668 43004
rect 2668 42948 2724 43004
rect 2724 42948 2728 43004
rect 2664 42944 2728 42948
rect 2744 43004 2808 43008
rect 2744 42948 2748 43004
rect 2748 42948 2804 43004
rect 2804 42948 2808 43004
rect 2744 42944 2808 42948
rect 2824 43004 2888 43008
rect 2824 42948 2828 43004
rect 2828 42948 2884 43004
rect 2884 42948 2888 43004
rect 2824 42944 2888 42948
rect 5847 43004 5911 43008
rect 5847 42948 5851 43004
rect 5851 42948 5907 43004
rect 5907 42948 5911 43004
rect 5847 42944 5911 42948
rect 5927 43004 5991 43008
rect 5927 42948 5931 43004
rect 5931 42948 5987 43004
rect 5987 42948 5991 43004
rect 5927 42944 5991 42948
rect 6007 43004 6071 43008
rect 6007 42948 6011 43004
rect 6011 42948 6067 43004
rect 6067 42948 6071 43004
rect 6007 42944 6071 42948
rect 6087 43004 6151 43008
rect 6087 42948 6091 43004
rect 6091 42948 6147 43004
rect 6147 42948 6151 43004
rect 6087 42944 6151 42948
rect 9111 43004 9175 43008
rect 9111 42948 9115 43004
rect 9115 42948 9171 43004
rect 9171 42948 9175 43004
rect 9111 42944 9175 42948
rect 9191 43004 9255 43008
rect 9191 42948 9195 43004
rect 9195 42948 9251 43004
rect 9251 42948 9255 43004
rect 9191 42944 9255 42948
rect 9271 43004 9335 43008
rect 9271 42948 9275 43004
rect 9275 42948 9331 43004
rect 9331 42948 9335 43004
rect 9271 42944 9335 42948
rect 9351 43004 9415 43008
rect 9351 42948 9355 43004
rect 9355 42948 9411 43004
rect 9411 42948 9415 43004
rect 9351 42944 9415 42948
rect 4215 42460 4279 42464
rect 4215 42404 4219 42460
rect 4219 42404 4275 42460
rect 4275 42404 4279 42460
rect 4215 42400 4279 42404
rect 4295 42460 4359 42464
rect 4295 42404 4299 42460
rect 4299 42404 4355 42460
rect 4355 42404 4359 42460
rect 4295 42400 4359 42404
rect 4375 42460 4439 42464
rect 4375 42404 4379 42460
rect 4379 42404 4435 42460
rect 4435 42404 4439 42460
rect 4375 42400 4439 42404
rect 4455 42460 4519 42464
rect 4455 42404 4459 42460
rect 4459 42404 4515 42460
rect 4515 42404 4519 42460
rect 4455 42400 4519 42404
rect 7479 42460 7543 42464
rect 7479 42404 7483 42460
rect 7483 42404 7539 42460
rect 7539 42404 7543 42460
rect 7479 42400 7543 42404
rect 7559 42460 7623 42464
rect 7559 42404 7563 42460
rect 7563 42404 7619 42460
rect 7619 42404 7623 42460
rect 7559 42400 7623 42404
rect 7639 42460 7703 42464
rect 7639 42404 7643 42460
rect 7643 42404 7699 42460
rect 7699 42404 7703 42460
rect 7639 42400 7703 42404
rect 7719 42460 7783 42464
rect 7719 42404 7723 42460
rect 7723 42404 7779 42460
rect 7779 42404 7783 42460
rect 7719 42400 7783 42404
rect 2584 41916 2648 41920
rect 2584 41860 2588 41916
rect 2588 41860 2644 41916
rect 2644 41860 2648 41916
rect 2584 41856 2648 41860
rect 2664 41916 2728 41920
rect 2664 41860 2668 41916
rect 2668 41860 2724 41916
rect 2724 41860 2728 41916
rect 2664 41856 2728 41860
rect 2744 41916 2808 41920
rect 2744 41860 2748 41916
rect 2748 41860 2804 41916
rect 2804 41860 2808 41916
rect 2744 41856 2808 41860
rect 2824 41916 2888 41920
rect 2824 41860 2828 41916
rect 2828 41860 2884 41916
rect 2884 41860 2888 41916
rect 2824 41856 2888 41860
rect 5847 41916 5911 41920
rect 5847 41860 5851 41916
rect 5851 41860 5907 41916
rect 5907 41860 5911 41916
rect 5847 41856 5911 41860
rect 5927 41916 5991 41920
rect 5927 41860 5931 41916
rect 5931 41860 5987 41916
rect 5987 41860 5991 41916
rect 5927 41856 5991 41860
rect 6007 41916 6071 41920
rect 6007 41860 6011 41916
rect 6011 41860 6067 41916
rect 6067 41860 6071 41916
rect 6007 41856 6071 41860
rect 6087 41916 6151 41920
rect 6087 41860 6091 41916
rect 6091 41860 6147 41916
rect 6147 41860 6151 41916
rect 6087 41856 6151 41860
rect 9111 41916 9175 41920
rect 9111 41860 9115 41916
rect 9115 41860 9171 41916
rect 9171 41860 9175 41916
rect 9111 41856 9175 41860
rect 9191 41916 9255 41920
rect 9191 41860 9195 41916
rect 9195 41860 9251 41916
rect 9251 41860 9255 41916
rect 9191 41856 9255 41860
rect 9271 41916 9335 41920
rect 9271 41860 9275 41916
rect 9275 41860 9331 41916
rect 9331 41860 9335 41916
rect 9271 41856 9335 41860
rect 9351 41916 9415 41920
rect 9351 41860 9355 41916
rect 9355 41860 9411 41916
rect 9411 41860 9415 41916
rect 9351 41856 9415 41860
rect 4660 41380 4724 41444
rect 4215 41372 4279 41376
rect 4215 41316 4219 41372
rect 4219 41316 4275 41372
rect 4275 41316 4279 41372
rect 4215 41312 4279 41316
rect 4295 41372 4359 41376
rect 4295 41316 4299 41372
rect 4299 41316 4355 41372
rect 4355 41316 4359 41372
rect 4295 41312 4359 41316
rect 4375 41372 4439 41376
rect 4375 41316 4379 41372
rect 4379 41316 4435 41372
rect 4435 41316 4439 41372
rect 4375 41312 4439 41316
rect 4455 41372 4519 41376
rect 4455 41316 4459 41372
rect 4459 41316 4515 41372
rect 4515 41316 4519 41372
rect 4455 41312 4519 41316
rect 7479 41372 7543 41376
rect 7479 41316 7483 41372
rect 7483 41316 7539 41372
rect 7539 41316 7543 41372
rect 7479 41312 7543 41316
rect 7559 41372 7623 41376
rect 7559 41316 7563 41372
rect 7563 41316 7619 41372
rect 7619 41316 7623 41372
rect 7559 41312 7623 41316
rect 7639 41372 7703 41376
rect 7639 41316 7643 41372
rect 7643 41316 7699 41372
rect 7699 41316 7703 41372
rect 7639 41312 7703 41316
rect 7719 41372 7783 41376
rect 7719 41316 7723 41372
rect 7723 41316 7779 41372
rect 7779 41316 7783 41372
rect 7719 41312 7783 41316
rect 2584 40828 2648 40832
rect 2584 40772 2588 40828
rect 2588 40772 2644 40828
rect 2644 40772 2648 40828
rect 2584 40768 2648 40772
rect 2664 40828 2728 40832
rect 2664 40772 2668 40828
rect 2668 40772 2724 40828
rect 2724 40772 2728 40828
rect 2664 40768 2728 40772
rect 2744 40828 2808 40832
rect 2744 40772 2748 40828
rect 2748 40772 2804 40828
rect 2804 40772 2808 40828
rect 2744 40768 2808 40772
rect 2824 40828 2888 40832
rect 2824 40772 2828 40828
rect 2828 40772 2884 40828
rect 2884 40772 2888 40828
rect 2824 40768 2888 40772
rect 5847 40828 5911 40832
rect 5847 40772 5851 40828
rect 5851 40772 5907 40828
rect 5907 40772 5911 40828
rect 5847 40768 5911 40772
rect 5927 40828 5991 40832
rect 5927 40772 5931 40828
rect 5931 40772 5987 40828
rect 5987 40772 5991 40828
rect 5927 40768 5991 40772
rect 6007 40828 6071 40832
rect 6007 40772 6011 40828
rect 6011 40772 6067 40828
rect 6067 40772 6071 40828
rect 6007 40768 6071 40772
rect 6087 40828 6151 40832
rect 6087 40772 6091 40828
rect 6091 40772 6147 40828
rect 6147 40772 6151 40828
rect 6087 40768 6151 40772
rect 9111 40828 9175 40832
rect 9111 40772 9115 40828
rect 9115 40772 9171 40828
rect 9171 40772 9175 40828
rect 9111 40768 9175 40772
rect 9191 40828 9255 40832
rect 9191 40772 9195 40828
rect 9195 40772 9251 40828
rect 9251 40772 9255 40828
rect 9191 40768 9255 40772
rect 9271 40828 9335 40832
rect 9271 40772 9275 40828
rect 9275 40772 9331 40828
rect 9331 40772 9335 40828
rect 9271 40768 9335 40772
rect 9351 40828 9415 40832
rect 9351 40772 9355 40828
rect 9355 40772 9411 40828
rect 9411 40772 9415 40828
rect 9351 40768 9415 40772
rect 2084 40292 2148 40356
rect 4215 40284 4279 40288
rect 4215 40228 4219 40284
rect 4219 40228 4275 40284
rect 4275 40228 4279 40284
rect 4215 40224 4279 40228
rect 4295 40284 4359 40288
rect 4295 40228 4299 40284
rect 4299 40228 4355 40284
rect 4355 40228 4359 40284
rect 4295 40224 4359 40228
rect 4375 40284 4439 40288
rect 4375 40228 4379 40284
rect 4379 40228 4435 40284
rect 4435 40228 4439 40284
rect 4375 40224 4439 40228
rect 4455 40284 4519 40288
rect 4455 40228 4459 40284
rect 4459 40228 4515 40284
rect 4515 40228 4519 40284
rect 4455 40224 4519 40228
rect 7479 40284 7543 40288
rect 7479 40228 7483 40284
rect 7483 40228 7539 40284
rect 7539 40228 7543 40284
rect 7479 40224 7543 40228
rect 7559 40284 7623 40288
rect 7559 40228 7563 40284
rect 7563 40228 7619 40284
rect 7619 40228 7623 40284
rect 7559 40224 7623 40228
rect 7639 40284 7703 40288
rect 7639 40228 7643 40284
rect 7643 40228 7699 40284
rect 7699 40228 7703 40284
rect 7639 40224 7703 40228
rect 7719 40284 7783 40288
rect 7719 40228 7723 40284
rect 7723 40228 7779 40284
rect 7779 40228 7783 40284
rect 7719 40224 7783 40228
rect 2268 40020 2332 40084
rect 2584 39740 2648 39744
rect 2584 39684 2588 39740
rect 2588 39684 2644 39740
rect 2644 39684 2648 39740
rect 2584 39680 2648 39684
rect 2664 39740 2728 39744
rect 2664 39684 2668 39740
rect 2668 39684 2724 39740
rect 2724 39684 2728 39740
rect 2664 39680 2728 39684
rect 2744 39740 2808 39744
rect 2744 39684 2748 39740
rect 2748 39684 2804 39740
rect 2804 39684 2808 39740
rect 2744 39680 2808 39684
rect 2824 39740 2888 39744
rect 2824 39684 2828 39740
rect 2828 39684 2884 39740
rect 2884 39684 2888 39740
rect 2824 39680 2888 39684
rect 5847 39740 5911 39744
rect 5847 39684 5851 39740
rect 5851 39684 5907 39740
rect 5907 39684 5911 39740
rect 5847 39680 5911 39684
rect 5927 39740 5991 39744
rect 5927 39684 5931 39740
rect 5931 39684 5987 39740
rect 5987 39684 5991 39740
rect 5927 39680 5991 39684
rect 6007 39740 6071 39744
rect 6007 39684 6011 39740
rect 6011 39684 6067 39740
rect 6067 39684 6071 39740
rect 6007 39680 6071 39684
rect 6087 39740 6151 39744
rect 6087 39684 6091 39740
rect 6091 39684 6147 39740
rect 6147 39684 6151 39740
rect 6087 39680 6151 39684
rect 9111 39740 9175 39744
rect 9111 39684 9115 39740
rect 9115 39684 9171 39740
rect 9171 39684 9175 39740
rect 9111 39680 9175 39684
rect 9191 39740 9255 39744
rect 9191 39684 9195 39740
rect 9195 39684 9251 39740
rect 9251 39684 9255 39740
rect 9191 39680 9255 39684
rect 9271 39740 9335 39744
rect 9271 39684 9275 39740
rect 9275 39684 9331 39740
rect 9331 39684 9335 39740
rect 9271 39680 9335 39684
rect 9351 39740 9415 39744
rect 9351 39684 9355 39740
rect 9355 39684 9411 39740
rect 9411 39684 9415 39740
rect 9351 39680 9415 39684
rect 4215 39196 4279 39200
rect 4215 39140 4219 39196
rect 4219 39140 4275 39196
rect 4275 39140 4279 39196
rect 4215 39136 4279 39140
rect 4295 39196 4359 39200
rect 4295 39140 4299 39196
rect 4299 39140 4355 39196
rect 4355 39140 4359 39196
rect 4295 39136 4359 39140
rect 4375 39196 4439 39200
rect 4375 39140 4379 39196
rect 4379 39140 4435 39196
rect 4435 39140 4439 39196
rect 4375 39136 4439 39140
rect 4455 39196 4519 39200
rect 4455 39140 4459 39196
rect 4459 39140 4515 39196
rect 4515 39140 4519 39196
rect 4455 39136 4519 39140
rect 7479 39196 7543 39200
rect 7479 39140 7483 39196
rect 7483 39140 7539 39196
rect 7539 39140 7543 39196
rect 7479 39136 7543 39140
rect 7559 39196 7623 39200
rect 7559 39140 7563 39196
rect 7563 39140 7619 39196
rect 7619 39140 7623 39196
rect 7559 39136 7623 39140
rect 7639 39196 7703 39200
rect 7639 39140 7643 39196
rect 7643 39140 7699 39196
rect 7699 39140 7703 39196
rect 7639 39136 7703 39140
rect 7719 39196 7783 39200
rect 7719 39140 7723 39196
rect 7723 39140 7779 39196
rect 7779 39140 7783 39196
rect 7719 39136 7783 39140
rect 2584 38652 2648 38656
rect 2584 38596 2588 38652
rect 2588 38596 2644 38652
rect 2644 38596 2648 38652
rect 2584 38592 2648 38596
rect 2664 38652 2728 38656
rect 2664 38596 2668 38652
rect 2668 38596 2724 38652
rect 2724 38596 2728 38652
rect 2664 38592 2728 38596
rect 2744 38652 2808 38656
rect 2744 38596 2748 38652
rect 2748 38596 2804 38652
rect 2804 38596 2808 38652
rect 2744 38592 2808 38596
rect 2824 38652 2888 38656
rect 2824 38596 2828 38652
rect 2828 38596 2884 38652
rect 2884 38596 2888 38652
rect 2824 38592 2888 38596
rect 5847 38652 5911 38656
rect 5847 38596 5851 38652
rect 5851 38596 5907 38652
rect 5907 38596 5911 38652
rect 5847 38592 5911 38596
rect 5927 38652 5991 38656
rect 5927 38596 5931 38652
rect 5931 38596 5987 38652
rect 5987 38596 5991 38652
rect 5927 38592 5991 38596
rect 6007 38652 6071 38656
rect 6007 38596 6011 38652
rect 6011 38596 6067 38652
rect 6067 38596 6071 38652
rect 6007 38592 6071 38596
rect 6087 38652 6151 38656
rect 6087 38596 6091 38652
rect 6091 38596 6147 38652
rect 6147 38596 6151 38652
rect 6087 38592 6151 38596
rect 9111 38652 9175 38656
rect 9111 38596 9115 38652
rect 9115 38596 9171 38652
rect 9171 38596 9175 38652
rect 9111 38592 9175 38596
rect 9191 38652 9255 38656
rect 9191 38596 9195 38652
rect 9195 38596 9251 38652
rect 9251 38596 9255 38652
rect 9191 38592 9255 38596
rect 9271 38652 9335 38656
rect 9271 38596 9275 38652
rect 9275 38596 9331 38652
rect 9331 38596 9335 38652
rect 9271 38592 9335 38596
rect 9351 38652 9415 38656
rect 9351 38596 9355 38652
rect 9355 38596 9411 38652
rect 9411 38596 9415 38652
rect 9351 38592 9415 38596
rect 4215 38108 4279 38112
rect 4215 38052 4219 38108
rect 4219 38052 4275 38108
rect 4275 38052 4279 38108
rect 4215 38048 4279 38052
rect 4295 38108 4359 38112
rect 4295 38052 4299 38108
rect 4299 38052 4355 38108
rect 4355 38052 4359 38108
rect 4295 38048 4359 38052
rect 4375 38108 4439 38112
rect 4375 38052 4379 38108
rect 4379 38052 4435 38108
rect 4435 38052 4439 38108
rect 4375 38048 4439 38052
rect 4455 38108 4519 38112
rect 4455 38052 4459 38108
rect 4459 38052 4515 38108
rect 4515 38052 4519 38108
rect 4455 38048 4519 38052
rect 7479 38108 7543 38112
rect 7479 38052 7483 38108
rect 7483 38052 7539 38108
rect 7539 38052 7543 38108
rect 7479 38048 7543 38052
rect 7559 38108 7623 38112
rect 7559 38052 7563 38108
rect 7563 38052 7619 38108
rect 7619 38052 7623 38108
rect 7559 38048 7623 38052
rect 7639 38108 7703 38112
rect 7639 38052 7643 38108
rect 7643 38052 7699 38108
rect 7699 38052 7703 38108
rect 7639 38048 7703 38052
rect 7719 38108 7783 38112
rect 7719 38052 7723 38108
rect 7723 38052 7779 38108
rect 7779 38052 7783 38108
rect 7719 38048 7783 38052
rect 2584 37564 2648 37568
rect 2584 37508 2588 37564
rect 2588 37508 2644 37564
rect 2644 37508 2648 37564
rect 2584 37504 2648 37508
rect 2664 37564 2728 37568
rect 2664 37508 2668 37564
rect 2668 37508 2724 37564
rect 2724 37508 2728 37564
rect 2664 37504 2728 37508
rect 2744 37564 2808 37568
rect 2744 37508 2748 37564
rect 2748 37508 2804 37564
rect 2804 37508 2808 37564
rect 2744 37504 2808 37508
rect 2824 37564 2888 37568
rect 2824 37508 2828 37564
rect 2828 37508 2884 37564
rect 2884 37508 2888 37564
rect 2824 37504 2888 37508
rect 5847 37564 5911 37568
rect 5847 37508 5851 37564
rect 5851 37508 5907 37564
rect 5907 37508 5911 37564
rect 5847 37504 5911 37508
rect 5927 37564 5991 37568
rect 5927 37508 5931 37564
rect 5931 37508 5987 37564
rect 5987 37508 5991 37564
rect 5927 37504 5991 37508
rect 6007 37564 6071 37568
rect 6007 37508 6011 37564
rect 6011 37508 6067 37564
rect 6067 37508 6071 37564
rect 6007 37504 6071 37508
rect 6087 37564 6151 37568
rect 6087 37508 6091 37564
rect 6091 37508 6147 37564
rect 6147 37508 6151 37564
rect 6087 37504 6151 37508
rect 9111 37564 9175 37568
rect 9111 37508 9115 37564
rect 9115 37508 9171 37564
rect 9171 37508 9175 37564
rect 9111 37504 9175 37508
rect 9191 37564 9255 37568
rect 9191 37508 9195 37564
rect 9195 37508 9251 37564
rect 9251 37508 9255 37564
rect 9191 37504 9255 37508
rect 9271 37564 9335 37568
rect 9271 37508 9275 37564
rect 9275 37508 9331 37564
rect 9331 37508 9335 37564
rect 9271 37504 9335 37508
rect 9351 37564 9415 37568
rect 9351 37508 9355 37564
rect 9355 37508 9411 37564
rect 9411 37508 9415 37564
rect 9351 37504 9415 37508
rect 4215 37020 4279 37024
rect 4215 36964 4219 37020
rect 4219 36964 4275 37020
rect 4275 36964 4279 37020
rect 4215 36960 4279 36964
rect 4295 37020 4359 37024
rect 4295 36964 4299 37020
rect 4299 36964 4355 37020
rect 4355 36964 4359 37020
rect 4295 36960 4359 36964
rect 4375 37020 4439 37024
rect 4375 36964 4379 37020
rect 4379 36964 4435 37020
rect 4435 36964 4439 37020
rect 4375 36960 4439 36964
rect 4455 37020 4519 37024
rect 4455 36964 4459 37020
rect 4459 36964 4515 37020
rect 4515 36964 4519 37020
rect 4455 36960 4519 36964
rect 7479 37020 7543 37024
rect 7479 36964 7483 37020
rect 7483 36964 7539 37020
rect 7539 36964 7543 37020
rect 7479 36960 7543 36964
rect 7559 37020 7623 37024
rect 7559 36964 7563 37020
rect 7563 36964 7619 37020
rect 7619 36964 7623 37020
rect 7559 36960 7623 36964
rect 7639 37020 7703 37024
rect 7639 36964 7643 37020
rect 7643 36964 7699 37020
rect 7699 36964 7703 37020
rect 7639 36960 7703 36964
rect 7719 37020 7783 37024
rect 7719 36964 7723 37020
rect 7723 36964 7779 37020
rect 7779 36964 7783 37020
rect 7719 36960 7783 36964
rect 2084 36756 2148 36820
rect 2584 36476 2648 36480
rect 2584 36420 2588 36476
rect 2588 36420 2644 36476
rect 2644 36420 2648 36476
rect 2584 36416 2648 36420
rect 2664 36476 2728 36480
rect 2664 36420 2668 36476
rect 2668 36420 2724 36476
rect 2724 36420 2728 36476
rect 2664 36416 2728 36420
rect 2744 36476 2808 36480
rect 2744 36420 2748 36476
rect 2748 36420 2804 36476
rect 2804 36420 2808 36476
rect 2744 36416 2808 36420
rect 2824 36476 2888 36480
rect 2824 36420 2828 36476
rect 2828 36420 2884 36476
rect 2884 36420 2888 36476
rect 2824 36416 2888 36420
rect 5847 36476 5911 36480
rect 5847 36420 5851 36476
rect 5851 36420 5907 36476
rect 5907 36420 5911 36476
rect 5847 36416 5911 36420
rect 5927 36476 5991 36480
rect 5927 36420 5931 36476
rect 5931 36420 5987 36476
rect 5987 36420 5991 36476
rect 5927 36416 5991 36420
rect 6007 36476 6071 36480
rect 6007 36420 6011 36476
rect 6011 36420 6067 36476
rect 6067 36420 6071 36476
rect 6007 36416 6071 36420
rect 6087 36476 6151 36480
rect 6087 36420 6091 36476
rect 6091 36420 6147 36476
rect 6147 36420 6151 36476
rect 6087 36416 6151 36420
rect 9111 36476 9175 36480
rect 9111 36420 9115 36476
rect 9115 36420 9171 36476
rect 9171 36420 9175 36476
rect 9111 36416 9175 36420
rect 9191 36476 9255 36480
rect 9191 36420 9195 36476
rect 9195 36420 9251 36476
rect 9251 36420 9255 36476
rect 9191 36416 9255 36420
rect 9271 36476 9335 36480
rect 9271 36420 9275 36476
rect 9275 36420 9331 36476
rect 9331 36420 9335 36476
rect 9271 36416 9335 36420
rect 9351 36476 9415 36480
rect 9351 36420 9355 36476
rect 9355 36420 9411 36476
rect 9411 36420 9415 36476
rect 9351 36416 9415 36420
rect 4215 35932 4279 35936
rect 4215 35876 4219 35932
rect 4219 35876 4275 35932
rect 4275 35876 4279 35932
rect 4215 35872 4279 35876
rect 4295 35932 4359 35936
rect 4295 35876 4299 35932
rect 4299 35876 4355 35932
rect 4355 35876 4359 35932
rect 4295 35872 4359 35876
rect 4375 35932 4439 35936
rect 4375 35876 4379 35932
rect 4379 35876 4435 35932
rect 4435 35876 4439 35932
rect 4375 35872 4439 35876
rect 4455 35932 4519 35936
rect 4455 35876 4459 35932
rect 4459 35876 4515 35932
rect 4515 35876 4519 35932
rect 4455 35872 4519 35876
rect 7479 35932 7543 35936
rect 7479 35876 7483 35932
rect 7483 35876 7539 35932
rect 7539 35876 7543 35932
rect 7479 35872 7543 35876
rect 7559 35932 7623 35936
rect 7559 35876 7563 35932
rect 7563 35876 7619 35932
rect 7619 35876 7623 35932
rect 7559 35872 7623 35876
rect 7639 35932 7703 35936
rect 7639 35876 7643 35932
rect 7643 35876 7699 35932
rect 7699 35876 7703 35932
rect 7639 35872 7703 35876
rect 7719 35932 7783 35936
rect 7719 35876 7723 35932
rect 7723 35876 7779 35932
rect 7779 35876 7783 35932
rect 7719 35872 7783 35876
rect 2584 35388 2648 35392
rect 2584 35332 2588 35388
rect 2588 35332 2644 35388
rect 2644 35332 2648 35388
rect 2584 35328 2648 35332
rect 2664 35388 2728 35392
rect 2664 35332 2668 35388
rect 2668 35332 2724 35388
rect 2724 35332 2728 35388
rect 2664 35328 2728 35332
rect 2744 35388 2808 35392
rect 2744 35332 2748 35388
rect 2748 35332 2804 35388
rect 2804 35332 2808 35388
rect 2744 35328 2808 35332
rect 2824 35388 2888 35392
rect 2824 35332 2828 35388
rect 2828 35332 2884 35388
rect 2884 35332 2888 35388
rect 2824 35328 2888 35332
rect 5847 35388 5911 35392
rect 5847 35332 5851 35388
rect 5851 35332 5907 35388
rect 5907 35332 5911 35388
rect 5847 35328 5911 35332
rect 5927 35388 5991 35392
rect 5927 35332 5931 35388
rect 5931 35332 5987 35388
rect 5987 35332 5991 35388
rect 5927 35328 5991 35332
rect 6007 35388 6071 35392
rect 6007 35332 6011 35388
rect 6011 35332 6067 35388
rect 6067 35332 6071 35388
rect 6007 35328 6071 35332
rect 6087 35388 6151 35392
rect 6087 35332 6091 35388
rect 6091 35332 6147 35388
rect 6147 35332 6151 35388
rect 6087 35328 6151 35332
rect 9111 35388 9175 35392
rect 9111 35332 9115 35388
rect 9115 35332 9171 35388
rect 9171 35332 9175 35388
rect 9111 35328 9175 35332
rect 9191 35388 9255 35392
rect 9191 35332 9195 35388
rect 9195 35332 9251 35388
rect 9251 35332 9255 35388
rect 9191 35328 9255 35332
rect 9271 35388 9335 35392
rect 9271 35332 9275 35388
rect 9275 35332 9331 35388
rect 9331 35332 9335 35388
rect 9271 35328 9335 35332
rect 9351 35388 9415 35392
rect 9351 35332 9355 35388
rect 9355 35332 9411 35388
rect 9411 35332 9415 35388
rect 9351 35328 9415 35332
rect 4215 34844 4279 34848
rect 4215 34788 4219 34844
rect 4219 34788 4275 34844
rect 4275 34788 4279 34844
rect 4215 34784 4279 34788
rect 4295 34844 4359 34848
rect 4295 34788 4299 34844
rect 4299 34788 4355 34844
rect 4355 34788 4359 34844
rect 4295 34784 4359 34788
rect 4375 34844 4439 34848
rect 4375 34788 4379 34844
rect 4379 34788 4435 34844
rect 4435 34788 4439 34844
rect 4375 34784 4439 34788
rect 4455 34844 4519 34848
rect 4455 34788 4459 34844
rect 4459 34788 4515 34844
rect 4515 34788 4519 34844
rect 4455 34784 4519 34788
rect 7479 34844 7543 34848
rect 7479 34788 7483 34844
rect 7483 34788 7539 34844
rect 7539 34788 7543 34844
rect 7479 34784 7543 34788
rect 7559 34844 7623 34848
rect 7559 34788 7563 34844
rect 7563 34788 7619 34844
rect 7619 34788 7623 34844
rect 7559 34784 7623 34788
rect 7639 34844 7703 34848
rect 7639 34788 7643 34844
rect 7643 34788 7699 34844
rect 7699 34788 7703 34844
rect 7639 34784 7703 34788
rect 7719 34844 7783 34848
rect 7719 34788 7723 34844
rect 7723 34788 7779 34844
rect 7779 34788 7783 34844
rect 7719 34784 7783 34788
rect 2584 34300 2648 34304
rect 2584 34244 2588 34300
rect 2588 34244 2644 34300
rect 2644 34244 2648 34300
rect 2584 34240 2648 34244
rect 2664 34300 2728 34304
rect 2664 34244 2668 34300
rect 2668 34244 2724 34300
rect 2724 34244 2728 34300
rect 2664 34240 2728 34244
rect 2744 34300 2808 34304
rect 2744 34244 2748 34300
rect 2748 34244 2804 34300
rect 2804 34244 2808 34300
rect 2744 34240 2808 34244
rect 2824 34300 2888 34304
rect 2824 34244 2828 34300
rect 2828 34244 2884 34300
rect 2884 34244 2888 34300
rect 2824 34240 2888 34244
rect 5847 34300 5911 34304
rect 5847 34244 5851 34300
rect 5851 34244 5907 34300
rect 5907 34244 5911 34300
rect 5847 34240 5911 34244
rect 5927 34300 5991 34304
rect 5927 34244 5931 34300
rect 5931 34244 5987 34300
rect 5987 34244 5991 34300
rect 5927 34240 5991 34244
rect 6007 34300 6071 34304
rect 6007 34244 6011 34300
rect 6011 34244 6067 34300
rect 6067 34244 6071 34300
rect 6007 34240 6071 34244
rect 6087 34300 6151 34304
rect 6087 34244 6091 34300
rect 6091 34244 6147 34300
rect 6147 34244 6151 34300
rect 6087 34240 6151 34244
rect 9111 34300 9175 34304
rect 9111 34244 9115 34300
rect 9115 34244 9171 34300
rect 9171 34244 9175 34300
rect 9111 34240 9175 34244
rect 9191 34300 9255 34304
rect 9191 34244 9195 34300
rect 9195 34244 9251 34300
rect 9251 34244 9255 34300
rect 9191 34240 9255 34244
rect 9271 34300 9335 34304
rect 9271 34244 9275 34300
rect 9275 34244 9331 34300
rect 9331 34244 9335 34300
rect 9271 34240 9335 34244
rect 9351 34300 9415 34304
rect 9351 34244 9355 34300
rect 9355 34244 9411 34300
rect 9411 34244 9415 34300
rect 9351 34240 9415 34244
rect 4215 33756 4279 33760
rect 4215 33700 4219 33756
rect 4219 33700 4275 33756
rect 4275 33700 4279 33756
rect 4215 33696 4279 33700
rect 4295 33756 4359 33760
rect 4295 33700 4299 33756
rect 4299 33700 4355 33756
rect 4355 33700 4359 33756
rect 4295 33696 4359 33700
rect 4375 33756 4439 33760
rect 4375 33700 4379 33756
rect 4379 33700 4435 33756
rect 4435 33700 4439 33756
rect 4375 33696 4439 33700
rect 4455 33756 4519 33760
rect 4455 33700 4459 33756
rect 4459 33700 4515 33756
rect 4515 33700 4519 33756
rect 4455 33696 4519 33700
rect 7479 33756 7543 33760
rect 7479 33700 7483 33756
rect 7483 33700 7539 33756
rect 7539 33700 7543 33756
rect 7479 33696 7543 33700
rect 7559 33756 7623 33760
rect 7559 33700 7563 33756
rect 7563 33700 7619 33756
rect 7619 33700 7623 33756
rect 7559 33696 7623 33700
rect 7639 33756 7703 33760
rect 7639 33700 7643 33756
rect 7643 33700 7699 33756
rect 7699 33700 7703 33756
rect 7639 33696 7703 33700
rect 7719 33756 7783 33760
rect 7719 33700 7723 33756
rect 7723 33700 7779 33756
rect 7779 33700 7783 33756
rect 7719 33696 7783 33700
rect 2584 33212 2648 33216
rect 2584 33156 2588 33212
rect 2588 33156 2644 33212
rect 2644 33156 2648 33212
rect 2584 33152 2648 33156
rect 2664 33212 2728 33216
rect 2664 33156 2668 33212
rect 2668 33156 2724 33212
rect 2724 33156 2728 33212
rect 2664 33152 2728 33156
rect 2744 33212 2808 33216
rect 2744 33156 2748 33212
rect 2748 33156 2804 33212
rect 2804 33156 2808 33212
rect 2744 33152 2808 33156
rect 2824 33212 2888 33216
rect 2824 33156 2828 33212
rect 2828 33156 2884 33212
rect 2884 33156 2888 33212
rect 2824 33152 2888 33156
rect 5847 33212 5911 33216
rect 5847 33156 5851 33212
rect 5851 33156 5907 33212
rect 5907 33156 5911 33212
rect 5847 33152 5911 33156
rect 5927 33212 5991 33216
rect 5927 33156 5931 33212
rect 5931 33156 5987 33212
rect 5987 33156 5991 33212
rect 5927 33152 5991 33156
rect 6007 33212 6071 33216
rect 6007 33156 6011 33212
rect 6011 33156 6067 33212
rect 6067 33156 6071 33212
rect 6007 33152 6071 33156
rect 6087 33212 6151 33216
rect 6087 33156 6091 33212
rect 6091 33156 6147 33212
rect 6147 33156 6151 33212
rect 6087 33152 6151 33156
rect 9111 33212 9175 33216
rect 9111 33156 9115 33212
rect 9115 33156 9171 33212
rect 9171 33156 9175 33212
rect 9111 33152 9175 33156
rect 9191 33212 9255 33216
rect 9191 33156 9195 33212
rect 9195 33156 9251 33212
rect 9251 33156 9255 33212
rect 9191 33152 9255 33156
rect 9271 33212 9335 33216
rect 9271 33156 9275 33212
rect 9275 33156 9331 33212
rect 9331 33156 9335 33212
rect 9271 33152 9335 33156
rect 9351 33212 9415 33216
rect 9351 33156 9355 33212
rect 9355 33156 9411 33212
rect 9411 33156 9415 33212
rect 9351 33152 9415 33156
rect 4215 32668 4279 32672
rect 4215 32612 4219 32668
rect 4219 32612 4275 32668
rect 4275 32612 4279 32668
rect 4215 32608 4279 32612
rect 4295 32668 4359 32672
rect 4295 32612 4299 32668
rect 4299 32612 4355 32668
rect 4355 32612 4359 32668
rect 4295 32608 4359 32612
rect 4375 32668 4439 32672
rect 4375 32612 4379 32668
rect 4379 32612 4435 32668
rect 4435 32612 4439 32668
rect 4375 32608 4439 32612
rect 4455 32668 4519 32672
rect 4455 32612 4459 32668
rect 4459 32612 4515 32668
rect 4515 32612 4519 32668
rect 4455 32608 4519 32612
rect 7479 32668 7543 32672
rect 7479 32612 7483 32668
rect 7483 32612 7539 32668
rect 7539 32612 7543 32668
rect 7479 32608 7543 32612
rect 7559 32668 7623 32672
rect 7559 32612 7563 32668
rect 7563 32612 7619 32668
rect 7619 32612 7623 32668
rect 7559 32608 7623 32612
rect 7639 32668 7703 32672
rect 7639 32612 7643 32668
rect 7643 32612 7699 32668
rect 7699 32612 7703 32668
rect 7639 32608 7703 32612
rect 7719 32668 7783 32672
rect 7719 32612 7723 32668
rect 7723 32612 7779 32668
rect 7779 32612 7783 32668
rect 7719 32608 7783 32612
rect 2584 32124 2648 32128
rect 2584 32068 2588 32124
rect 2588 32068 2644 32124
rect 2644 32068 2648 32124
rect 2584 32064 2648 32068
rect 2664 32124 2728 32128
rect 2664 32068 2668 32124
rect 2668 32068 2724 32124
rect 2724 32068 2728 32124
rect 2664 32064 2728 32068
rect 2744 32124 2808 32128
rect 2744 32068 2748 32124
rect 2748 32068 2804 32124
rect 2804 32068 2808 32124
rect 2744 32064 2808 32068
rect 2824 32124 2888 32128
rect 2824 32068 2828 32124
rect 2828 32068 2884 32124
rect 2884 32068 2888 32124
rect 2824 32064 2888 32068
rect 5847 32124 5911 32128
rect 5847 32068 5851 32124
rect 5851 32068 5907 32124
rect 5907 32068 5911 32124
rect 5847 32064 5911 32068
rect 5927 32124 5991 32128
rect 5927 32068 5931 32124
rect 5931 32068 5987 32124
rect 5987 32068 5991 32124
rect 5927 32064 5991 32068
rect 6007 32124 6071 32128
rect 6007 32068 6011 32124
rect 6011 32068 6067 32124
rect 6067 32068 6071 32124
rect 6007 32064 6071 32068
rect 6087 32124 6151 32128
rect 6087 32068 6091 32124
rect 6091 32068 6147 32124
rect 6147 32068 6151 32124
rect 6087 32064 6151 32068
rect 9111 32124 9175 32128
rect 9111 32068 9115 32124
rect 9115 32068 9171 32124
rect 9171 32068 9175 32124
rect 9111 32064 9175 32068
rect 9191 32124 9255 32128
rect 9191 32068 9195 32124
rect 9195 32068 9251 32124
rect 9251 32068 9255 32124
rect 9191 32064 9255 32068
rect 9271 32124 9335 32128
rect 9271 32068 9275 32124
rect 9275 32068 9331 32124
rect 9331 32068 9335 32124
rect 9271 32064 9335 32068
rect 9351 32124 9415 32128
rect 9351 32068 9355 32124
rect 9355 32068 9411 32124
rect 9411 32068 9415 32124
rect 9351 32064 9415 32068
rect 4215 31580 4279 31584
rect 4215 31524 4219 31580
rect 4219 31524 4275 31580
rect 4275 31524 4279 31580
rect 4215 31520 4279 31524
rect 4295 31580 4359 31584
rect 4295 31524 4299 31580
rect 4299 31524 4355 31580
rect 4355 31524 4359 31580
rect 4295 31520 4359 31524
rect 4375 31580 4439 31584
rect 4375 31524 4379 31580
rect 4379 31524 4435 31580
rect 4435 31524 4439 31580
rect 4375 31520 4439 31524
rect 4455 31580 4519 31584
rect 4455 31524 4459 31580
rect 4459 31524 4515 31580
rect 4515 31524 4519 31580
rect 4455 31520 4519 31524
rect 7479 31580 7543 31584
rect 7479 31524 7483 31580
rect 7483 31524 7539 31580
rect 7539 31524 7543 31580
rect 7479 31520 7543 31524
rect 7559 31580 7623 31584
rect 7559 31524 7563 31580
rect 7563 31524 7619 31580
rect 7619 31524 7623 31580
rect 7559 31520 7623 31524
rect 7639 31580 7703 31584
rect 7639 31524 7643 31580
rect 7643 31524 7699 31580
rect 7699 31524 7703 31580
rect 7639 31520 7703 31524
rect 7719 31580 7783 31584
rect 7719 31524 7723 31580
rect 7723 31524 7779 31580
rect 7779 31524 7783 31580
rect 7719 31520 7783 31524
rect 2584 31036 2648 31040
rect 2584 30980 2588 31036
rect 2588 30980 2644 31036
rect 2644 30980 2648 31036
rect 2584 30976 2648 30980
rect 2664 31036 2728 31040
rect 2664 30980 2668 31036
rect 2668 30980 2724 31036
rect 2724 30980 2728 31036
rect 2664 30976 2728 30980
rect 2744 31036 2808 31040
rect 2744 30980 2748 31036
rect 2748 30980 2804 31036
rect 2804 30980 2808 31036
rect 2744 30976 2808 30980
rect 2824 31036 2888 31040
rect 2824 30980 2828 31036
rect 2828 30980 2884 31036
rect 2884 30980 2888 31036
rect 2824 30976 2888 30980
rect 5847 31036 5911 31040
rect 5847 30980 5851 31036
rect 5851 30980 5907 31036
rect 5907 30980 5911 31036
rect 5847 30976 5911 30980
rect 5927 31036 5991 31040
rect 5927 30980 5931 31036
rect 5931 30980 5987 31036
rect 5987 30980 5991 31036
rect 5927 30976 5991 30980
rect 6007 31036 6071 31040
rect 6007 30980 6011 31036
rect 6011 30980 6067 31036
rect 6067 30980 6071 31036
rect 6007 30976 6071 30980
rect 6087 31036 6151 31040
rect 6087 30980 6091 31036
rect 6091 30980 6147 31036
rect 6147 30980 6151 31036
rect 6087 30976 6151 30980
rect 9111 31036 9175 31040
rect 9111 30980 9115 31036
rect 9115 30980 9171 31036
rect 9171 30980 9175 31036
rect 9111 30976 9175 30980
rect 9191 31036 9255 31040
rect 9191 30980 9195 31036
rect 9195 30980 9251 31036
rect 9251 30980 9255 31036
rect 9191 30976 9255 30980
rect 9271 31036 9335 31040
rect 9271 30980 9275 31036
rect 9275 30980 9331 31036
rect 9331 30980 9335 31036
rect 9271 30976 9335 30980
rect 9351 31036 9415 31040
rect 9351 30980 9355 31036
rect 9355 30980 9411 31036
rect 9411 30980 9415 31036
rect 9351 30976 9415 30980
rect 4215 30492 4279 30496
rect 4215 30436 4219 30492
rect 4219 30436 4275 30492
rect 4275 30436 4279 30492
rect 4215 30432 4279 30436
rect 4295 30492 4359 30496
rect 4295 30436 4299 30492
rect 4299 30436 4355 30492
rect 4355 30436 4359 30492
rect 4295 30432 4359 30436
rect 4375 30492 4439 30496
rect 4375 30436 4379 30492
rect 4379 30436 4435 30492
rect 4435 30436 4439 30492
rect 4375 30432 4439 30436
rect 4455 30492 4519 30496
rect 4455 30436 4459 30492
rect 4459 30436 4515 30492
rect 4515 30436 4519 30492
rect 4455 30432 4519 30436
rect 7479 30492 7543 30496
rect 7479 30436 7483 30492
rect 7483 30436 7539 30492
rect 7539 30436 7543 30492
rect 7479 30432 7543 30436
rect 7559 30492 7623 30496
rect 7559 30436 7563 30492
rect 7563 30436 7619 30492
rect 7619 30436 7623 30492
rect 7559 30432 7623 30436
rect 7639 30492 7703 30496
rect 7639 30436 7643 30492
rect 7643 30436 7699 30492
rect 7699 30436 7703 30492
rect 7639 30432 7703 30436
rect 7719 30492 7783 30496
rect 7719 30436 7723 30492
rect 7723 30436 7779 30492
rect 7779 30436 7783 30492
rect 7719 30432 7783 30436
rect 2584 29948 2648 29952
rect 2584 29892 2588 29948
rect 2588 29892 2644 29948
rect 2644 29892 2648 29948
rect 2584 29888 2648 29892
rect 2664 29948 2728 29952
rect 2664 29892 2668 29948
rect 2668 29892 2724 29948
rect 2724 29892 2728 29948
rect 2664 29888 2728 29892
rect 2744 29948 2808 29952
rect 2744 29892 2748 29948
rect 2748 29892 2804 29948
rect 2804 29892 2808 29948
rect 2744 29888 2808 29892
rect 2824 29948 2888 29952
rect 2824 29892 2828 29948
rect 2828 29892 2884 29948
rect 2884 29892 2888 29948
rect 2824 29888 2888 29892
rect 5847 29948 5911 29952
rect 5847 29892 5851 29948
rect 5851 29892 5907 29948
rect 5907 29892 5911 29948
rect 5847 29888 5911 29892
rect 5927 29948 5991 29952
rect 5927 29892 5931 29948
rect 5931 29892 5987 29948
rect 5987 29892 5991 29948
rect 5927 29888 5991 29892
rect 6007 29948 6071 29952
rect 6007 29892 6011 29948
rect 6011 29892 6067 29948
rect 6067 29892 6071 29948
rect 6007 29888 6071 29892
rect 6087 29948 6151 29952
rect 6087 29892 6091 29948
rect 6091 29892 6147 29948
rect 6147 29892 6151 29948
rect 6087 29888 6151 29892
rect 9111 29948 9175 29952
rect 9111 29892 9115 29948
rect 9115 29892 9171 29948
rect 9171 29892 9175 29948
rect 9111 29888 9175 29892
rect 9191 29948 9255 29952
rect 9191 29892 9195 29948
rect 9195 29892 9251 29948
rect 9251 29892 9255 29948
rect 9191 29888 9255 29892
rect 9271 29948 9335 29952
rect 9271 29892 9275 29948
rect 9275 29892 9331 29948
rect 9331 29892 9335 29948
rect 9271 29888 9335 29892
rect 9351 29948 9415 29952
rect 9351 29892 9355 29948
rect 9355 29892 9411 29948
rect 9411 29892 9415 29948
rect 9351 29888 9415 29892
rect 4215 29404 4279 29408
rect 4215 29348 4219 29404
rect 4219 29348 4275 29404
rect 4275 29348 4279 29404
rect 4215 29344 4279 29348
rect 4295 29404 4359 29408
rect 4295 29348 4299 29404
rect 4299 29348 4355 29404
rect 4355 29348 4359 29404
rect 4295 29344 4359 29348
rect 4375 29404 4439 29408
rect 4375 29348 4379 29404
rect 4379 29348 4435 29404
rect 4435 29348 4439 29404
rect 4375 29344 4439 29348
rect 4455 29404 4519 29408
rect 4455 29348 4459 29404
rect 4459 29348 4515 29404
rect 4515 29348 4519 29404
rect 4455 29344 4519 29348
rect 7479 29404 7543 29408
rect 7479 29348 7483 29404
rect 7483 29348 7539 29404
rect 7539 29348 7543 29404
rect 7479 29344 7543 29348
rect 7559 29404 7623 29408
rect 7559 29348 7563 29404
rect 7563 29348 7619 29404
rect 7619 29348 7623 29404
rect 7559 29344 7623 29348
rect 7639 29404 7703 29408
rect 7639 29348 7643 29404
rect 7643 29348 7699 29404
rect 7699 29348 7703 29404
rect 7639 29344 7703 29348
rect 7719 29404 7783 29408
rect 7719 29348 7723 29404
rect 7723 29348 7779 29404
rect 7779 29348 7783 29404
rect 7719 29344 7783 29348
rect 2584 28860 2648 28864
rect 2584 28804 2588 28860
rect 2588 28804 2644 28860
rect 2644 28804 2648 28860
rect 2584 28800 2648 28804
rect 2664 28860 2728 28864
rect 2664 28804 2668 28860
rect 2668 28804 2724 28860
rect 2724 28804 2728 28860
rect 2664 28800 2728 28804
rect 2744 28860 2808 28864
rect 2744 28804 2748 28860
rect 2748 28804 2804 28860
rect 2804 28804 2808 28860
rect 2744 28800 2808 28804
rect 2824 28860 2888 28864
rect 2824 28804 2828 28860
rect 2828 28804 2884 28860
rect 2884 28804 2888 28860
rect 2824 28800 2888 28804
rect 5847 28860 5911 28864
rect 5847 28804 5851 28860
rect 5851 28804 5907 28860
rect 5907 28804 5911 28860
rect 5847 28800 5911 28804
rect 5927 28860 5991 28864
rect 5927 28804 5931 28860
rect 5931 28804 5987 28860
rect 5987 28804 5991 28860
rect 5927 28800 5991 28804
rect 6007 28860 6071 28864
rect 6007 28804 6011 28860
rect 6011 28804 6067 28860
rect 6067 28804 6071 28860
rect 6007 28800 6071 28804
rect 6087 28860 6151 28864
rect 6087 28804 6091 28860
rect 6091 28804 6147 28860
rect 6147 28804 6151 28860
rect 6087 28800 6151 28804
rect 9111 28860 9175 28864
rect 9111 28804 9115 28860
rect 9115 28804 9171 28860
rect 9171 28804 9175 28860
rect 9111 28800 9175 28804
rect 9191 28860 9255 28864
rect 9191 28804 9195 28860
rect 9195 28804 9251 28860
rect 9251 28804 9255 28860
rect 9191 28800 9255 28804
rect 9271 28860 9335 28864
rect 9271 28804 9275 28860
rect 9275 28804 9331 28860
rect 9331 28804 9335 28860
rect 9271 28800 9335 28804
rect 9351 28860 9415 28864
rect 9351 28804 9355 28860
rect 9355 28804 9411 28860
rect 9411 28804 9415 28860
rect 9351 28800 9415 28804
rect 4215 28316 4279 28320
rect 4215 28260 4219 28316
rect 4219 28260 4275 28316
rect 4275 28260 4279 28316
rect 4215 28256 4279 28260
rect 4295 28316 4359 28320
rect 4295 28260 4299 28316
rect 4299 28260 4355 28316
rect 4355 28260 4359 28316
rect 4295 28256 4359 28260
rect 4375 28316 4439 28320
rect 4375 28260 4379 28316
rect 4379 28260 4435 28316
rect 4435 28260 4439 28316
rect 4375 28256 4439 28260
rect 4455 28316 4519 28320
rect 4455 28260 4459 28316
rect 4459 28260 4515 28316
rect 4515 28260 4519 28316
rect 4455 28256 4519 28260
rect 7479 28316 7543 28320
rect 7479 28260 7483 28316
rect 7483 28260 7539 28316
rect 7539 28260 7543 28316
rect 7479 28256 7543 28260
rect 7559 28316 7623 28320
rect 7559 28260 7563 28316
rect 7563 28260 7619 28316
rect 7619 28260 7623 28316
rect 7559 28256 7623 28260
rect 7639 28316 7703 28320
rect 7639 28260 7643 28316
rect 7643 28260 7699 28316
rect 7699 28260 7703 28316
rect 7639 28256 7703 28260
rect 7719 28316 7783 28320
rect 7719 28260 7723 28316
rect 7723 28260 7779 28316
rect 7779 28260 7783 28316
rect 7719 28256 7783 28260
rect 2584 27772 2648 27776
rect 2584 27716 2588 27772
rect 2588 27716 2644 27772
rect 2644 27716 2648 27772
rect 2584 27712 2648 27716
rect 2664 27772 2728 27776
rect 2664 27716 2668 27772
rect 2668 27716 2724 27772
rect 2724 27716 2728 27772
rect 2664 27712 2728 27716
rect 2744 27772 2808 27776
rect 2744 27716 2748 27772
rect 2748 27716 2804 27772
rect 2804 27716 2808 27772
rect 2744 27712 2808 27716
rect 2824 27772 2888 27776
rect 2824 27716 2828 27772
rect 2828 27716 2884 27772
rect 2884 27716 2888 27772
rect 2824 27712 2888 27716
rect 5847 27772 5911 27776
rect 5847 27716 5851 27772
rect 5851 27716 5907 27772
rect 5907 27716 5911 27772
rect 5847 27712 5911 27716
rect 5927 27772 5991 27776
rect 5927 27716 5931 27772
rect 5931 27716 5987 27772
rect 5987 27716 5991 27772
rect 5927 27712 5991 27716
rect 6007 27772 6071 27776
rect 6007 27716 6011 27772
rect 6011 27716 6067 27772
rect 6067 27716 6071 27772
rect 6007 27712 6071 27716
rect 6087 27772 6151 27776
rect 6087 27716 6091 27772
rect 6091 27716 6147 27772
rect 6147 27716 6151 27772
rect 6087 27712 6151 27716
rect 9111 27772 9175 27776
rect 9111 27716 9115 27772
rect 9115 27716 9171 27772
rect 9171 27716 9175 27772
rect 9111 27712 9175 27716
rect 9191 27772 9255 27776
rect 9191 27716 9195 27772
rect 9195 27716 9251 27772
rect 9251 27716 9255 27772
rect 9191 27712 9255 27716
rect 9271 27772 9335 27776
rect 9271 27716 9275 27772
rect 9275 27716 9331 27772
rect 9331 27716 9335 27772
rect 9271 27712 9335 27716
rect 9351 27772 9415 27776
rect 9351 27716 9355 27772
rect 9355 27716 9411 27772
rect 9411 27716 9415 27772
rect 9351 27712 9415 27716
rect 4215 27228 4279 27232
rect 4215 27172 4219 27228
rect 4219 27172 4275 27228
rect 4275 27172 4279 27228
rect 4215 27168 4279 27172
rect 4295 27228 4359 27232
rect 4295 27172 4299 27228
rect 4299 27172 4355 27228
rect 4355 27172 4359 27228
rect 4295 27168 4359 27172
rect 4375 27228 4439 27232
rect 4375 27172 4379 27228
rect 4379 27172 4435 27228
rect 4435 27172 4439 27228
rect 4375 27168 4439 27172
rect 4455 27228 4519 27232
rect 4455 27172 4459 27228
rect 4459 27172 4515 27228
rect 4515 27172 4519 27228
rect 4455 27168 4519 27172
rect 7479 27228 7543 27232
rect 7479 27172 7483 27228
rect 7483 27172 7539 27228
rect 7539 27172 7543 27228
rect 7479 27168 7543 27172
rect 7559 27228 7623 27232
rect 7559 27172 7563 27228
rect 7563 27172 7619 27228
rect 7619 27172 7623 27228
rect 7559 27168 7623 27172
rect 7639 27228 7703 27232
rect 7639 27172 7643 27228
rect 7643 27172 7699 27228
rect 7699 27172 7703 27228
rect 7639 27168 7703 27172
rect 7719 27228 7783 27232
rect 7719 27172 7723 27228
rect 7723 27172 7779 27228
rect 7779 27172 7783 27228
rect 7719 27168 7783 27172
rect 2584 26684 2648 26688
rect 2584 26628 2588 26684
rect 2588 26628 2644 26684
rect 2644 26628 2648 26684
rect 2584 26624 2648 26628
rect 2664 26684 2728 26688
rect 2664 26628 2668 26684
rect 2668 26628 2724 26684
rect 2724 26628 2728 26684
rect 2664 26624 2728 26628
rect 2744 26684 2808 26688
rect 2744 26628 2748 26684
rect 2748 26628 2804 26684
rect 2804 26628 2808 26684
rect 2744 26624 2808 26628
rect 2824 26684 2888 26688
rect 2824 26628 2828 26684
rect 2828 26628 2884 26684
rect 2884 26628 2888 26684
rect 2824 26624 2888 26628
rect 5847 26684 5911 26688
rect 5847 26628 5851 26684
rect 5851 26628 5907 26684
rect 5907 26628 5911 26684
rect 5847 26624 5911 26628
rect 5927 26684 5991 26688
rect 5927 26628 5931 26684
rect 5931 26628 5987 26684
rect 5987 26628 5991 26684
rect 5927 26624 5991 26628
rect 6007 26684 6071 26688
rect 6007 26628 6011 26684
rect 6011 26628 6067 26684
rect 6067 26628 6071 26684
rect 6007 26624 6071 26628
rect 6087 26684 6151 26688
rect 6087 26628 6091 26684
rect 6091 26628 6147 26684
rect 6147 26628 6151 26684
rect 6087 26624 6151 26628
rect 9111 26684 9175 26688
rect 9111 26628 9115 26684
rect 9115 26628 9171 26684
rect 9171 26628 9175 26684
rect 9111 26624 9175 26628
rect 9191 26684 9255 26688
rect 9191 26628 9195 26684
rect 9195 26628 9251 26684
rect 9251 26628 9255 26684
rect 9191 26624 9255 26628
rect 9271 26684 9335 26688
rect 9271 26628 9275 26684
rect 9275 26628 9331 26684
rect 9331 26628 9335 26684
rect 9271 26624 9335 26628
rect 9351 26684 9415 26688
rect 9351 26628 9355 26684
rect 9355 26628 9411 26684
rect 9411 26628 9415 26684
rect 9351 26624 9415 26628
rect 4215 26140 4279 26144
rect 4215 26084 4219 26140
rect 4219 26084 4275 26140
rect 4275 26084 4279 26140
rect 4215 26080 4279 26084
rect 4295 26140 4359 26144
rect 4295 26084 4299 26140
rect 4299 26084 4355 26140
rect 4355 26084 4359 26140
rect 4295 26080 4359 26084
rect 4375 26140 4439 26144
rect 4375 26084 4379 26140
rect 4379 26084 4435 26140
rect 4435 26084 4439 26140
rect 4375 26080 4439 26084
rect 4455 26140 4519 26144
rect 4455 26084 4459 26140
rect 4459 26084 4515 26140
rect 4515 26084 4519 26140
rect 4455 26080 4519 26084
rect 7479 26140 7543 26144
rect 7479 26084 7483 26140
rect 7483 26084 7539 26140
rect 7539 26084 7543 26140
rect 7479 26080 7543 26084
rect 7559 26140 7623 26144
rect 7559 26084 7563 26140
rect 7563 26084 7619 26140
rect 7619 26084 7623 26140
rect 7559 26080 7623 26084
rect 7639 26140 7703 26144
rect 7639 26084 7643 26140
rect 7643 26084 7699 26140
rect 7699 26084 7703 26140
rect 7639 26080 7703 26084
rect 7719 26140 7783 26144
rect 7719 26084 7723 26140
rect 7723 26084 7779 26140
rect 7779 26084 7783 26140
rect 7719 26080 7783 26084
rect 2584 25596 2648 25600
rect 2584 25540 2588 25596
rect 2588 25540 2644 25596
rect 2644 25540 2648 25596
rect 2584 25536 2648 25540
rect 2664 25596 2728 25600
rect 2664 25540 2668 25596
rect 2668 25540 2724 25596
rect 2724 25540 2728 25596
rect 2664 25536 2728 25540
rect 2744 25596 2808 25600
rect 2744 25540 2748 25596
rect 2748 25540 2804 25596
rect 2804 25540 2808 25596
rect 2744 25536 2808 25540
rect 2824 25596 2888 25600
rect 2824 25540 2828 25596
rect 2828 25540 2884 25596
rect 2884 25540 2888 25596
rect 2824 25536 2888 25540
rect 5847 25596 5911 25600
rect 5847 25540 5851 25596
rect 5851 25540 5907 25596
rect 5907 25540 5911 25596
rect 5847 25536 5911 25540
rect 5927 25596 5991 25600
rect 5927 25540 5931 25596
rect 5931 25540 5987 25596
rect 5987 25540 5991 25596
rect 5927 25536 5991 25540
rect 6007 25596 6071 25600
rect 6007 25540 6011 25596
rect 6011 25540 6067 25596
rect 6067 25540 6071 25596
rect 6007 25536 6071 25540
rect 6087 25596 6151 25600
rect 6087 25540 6091 25596
rect 6091 25540 6147 25596
rect 6147 25540 6151 25596
rect 6087 25536 6151 25540
rect 9111 25596 9175 25600
rect 9111 25540 9115 25596
rect 9115 25540 9171 25596
rect 9171 25540 9175 25596
rect 9111 25536 9175 25540
rect 9191 25596 9255 25600
rect 9191 25540 9195 25596
rect 9195 25540 9251 25596
rect 9251 25540 9255 25596
rect 9191 25536 9255 25540
rect 9271 25596 9335 25600
rect 9271 25540 9275 25596
rect 9275 25540 9331 25596
rect 9331 25540 9335 25596
rect 9271 25536 9335 25540
rect 9351 25596 9415 25600
rect 9351 25540 9355 25596
rect 9355 25540 9411 25596
rect 9411 25540 9415 25596
rect 9351 25536 9415 25540
rect 4215 25052 4279 25056
rect 4215 24996 4219 25052
rect 4219 24996 4275 25052
rect 4275 24996 4279 25052
rect 4215 24992 4279 24996
rect 4295 25052 4359 25056
rect 4295 24996 4299 25052
rect 4299 24996 4355 25052
rect 4355 24996 4359 25052
rect 4295 24992 4359 24996
rect 4375 25052 4439 25056
rect 4375 24996 4379 25052
rect 4379 24996 4435 25052
rect 4435 24996 4439 25052
rect 4375 24992 4439 24996
rect 4455 25052 4519 25056
rect 4455 24996 4459 25052
rect 4459 24996 4515 25052
rect 4515 24996 4519 25052
rect 4455 24992 4519 24996
rect 7479 25052 7543 25056
rect 7479 24996 7483 25052
rect 7483 24996 7539 25052
rect 7539 24996 7543 25052
rect 7479 24992 7543 24996
rect 7559 25052 7623 25056
rect 7559 24996 7563 25052
rect 7563 24996 7619 25052
rect 7619 24996 7623 25052
rect 7559 24992 7623 24996
rect 7639 25052 7703 25056
rect 7639 24996 7643 25052
rect 7643 24996 7699 25052
rect 7699 24996 7703 25052
rect 7639 24992 7703 24996
rect 7719 25052 7783 25056
rect 7719 24996 7723 25052
rect 7723 24996 7779 25052
rect 7779 24996 7783 25052
rect 7719 24992 7783 24996
rect 2584 24508 2648 24512
rect 2584 24452 2588 24508
rect 2588 24452 2644 24508
rect 2644 24452 2648 24508
rect 2584 24448 2648 24452
rect 2664 24508 2728 24512
rect 2664 24452 2668 24508
rect 2668 24452 2724 24508
rect 2724 24452 2728 24508
rect 2664 24448 2728 24452
rect 2744 24508 2808 24512
rect 2744 24452 2748 24508
rect 2748 24452 2804 24508
rect 2804 24452 2808 24508
rect 2744 24448 2808 24452
rect 2824 24508 2888 24512
rect 2824 24452 2828 24508
rect 2828 24452 2884 24508
rect 2884 24452 2888 24508
rect 2824 24448 2888 24452
rect 5847 24508 5911 24512
rect 5847 24452 5851 24508
rect 5851 24452 5907 24508
rect 5907 24452 5911 24508
rect 5847 24448 5911 24452
rect 5927 24508 5991 24512
rect 5927 24452 5931 24508
rect 5931 24452 5987 24508
rect 5987 24452 5991 24508
rect 5927 24448 5991 24452
rect 6007 24508 6071 24512
rect 6007 24452 6011 24508
rect 6011 24452 6067 24508
rect 6067 24452 6071 24508
rect 6007 24448 6071 24452
rect 6087 24508 6151 24512
rect 6087 24452 6091 24508
rect 6091 24452 6147 24508
rect 6147 24452 6151 24508
rect 6087 24448 6151 24452
rect 9111 24508 9175 24512
rect 9111 24452 9115 24508
rect 9115 24452 9171 24508
rect 9171 24452 9175 24508
rect 9111 24448 9175 24452
rect 9191 24508 9255 24512
rect 9191 24452 9195 24508
rect 9195 24452 9251 24508
rect 9251 24452 9255 24508
rect 9191 24448 9255 24452
rect 9271 24508 9335 24512
rect 9271 24452 9275 24508
rect 9275 24452 9331 24508
rect 9331 24452 9335 24508
rect 9271 24448 9335 24452
rect 9351 24508 9415 24512
rect 9351 24452 9355 24508
rect 9355 24452 9411 24508
rect 9411 24452 9415 24508
rect 9351 24448 9415 24452
rect 4215 23964 4279 23968
rect 4215 23908 4219 23964
rect 4219 23908 4275 23964
rect 4275 23908 4279 23964
rect 4215 23904 4279 23908
rect 4295 23964 4359 23968
rect 4295 23908 4299 23964
rect 4299 23908 4355 23964
rect 4355 23908 4359 23964
rect 4295 23904 4359 23908
rect 4375 23964 4439 23968
rect 4375 23908 4379 23964
rect 4379 23908 4435 23964
rect 4435 23908 4439 23964
rect 4375 23904 4439 23908
rect 4455 23964 4519 23968
rect 4455 23908 4459 23964
rect 4459 23908 4515 23964
rect 4515 23908 4519 23964
rect 4455 23904 4519 23908
rect 7479 23964 7543 23968
rect 7479 23908 7483 23964
rect 7483 23908 7539 23964
rect 7539 23908 7543 23964
rect 7479 23904 7543 23908
rect 7559 23964 7623 23968
rect 7559 23908 7563 23964
rect 7563 23908 7619 23964
rect 7619 23908 7623 23964
rect 7559 23904 7623 23908
rect 7639 23964 7703 23968
rect 7639 23908 7643 23964
rect 7643 23908 7699 23964
rect 7699 23908 7703 23964
rect 7639 23904 7703 23908
rect 7719 23964 7783 23968
rect 7719 23908 7723 23964
rect 7723 23908 7779 23964
rect 7779 23908 7783 23964
rect 7719 23904 7783 23908
rect 1164 23564 1228 23628
rect 2584 23420 2648 23424
rect 2584 23364 2588 23420
rect 2588 23364 2644 23420
rect 2644 23364 2648 23420
rect 2584 23360 2648 23364
rect 2664 23420 2728 23424
rect 2664 23364 2668 23420
rect 2668 23364 2724 23420
rect 2724 23364 2728 23420
rect 2664 23360 2728 23364
rect 2744 23420 2808 23424
rect 2744 23364 2748 23420
rect 2748 23364 2804 23420
rect 2804 23364 2808 23420
rect 2744 23360 2808 23364
rect 2824 23420 2888 23424
rect 2824 23364 2828 23420
rect 2828 23364 2884 23420
rect 2884 23364 2888 23420
rect 2824 23360 2888 23364
rect 5847 23420 5911 23424
rect 5847 23364 5851 23420
rect 5851 23364 5907 23420
rect 5907 23364 5911 23420
rect 5847 23360 5911 23364
rect 5927 23420 5991 23424
rect 5927 23364 5931 23420
rect 5931 23364 5987 23420
rect 5987 23364 5991 23420
rect 5927 23360 5991 23364
rect 6007 23420 6071 23424
rect 6007 23364 6011 23420
rect 6011 23364 6067 23420
rect 6067 23364 6071 23420
rect 6007 23360 6071 23364
rect 6087 23420 6151 23424
rect 6087 23364 6091 23420
rect 6091 23364 6147 23420
rect 6147 23364 6151 23420
rect 6087 23360 6151 23364
rect 9111 23420 9175 23424
rect 9111 23364 9115 23420
rect 9115 23364 9171 23420
rect 9171 23364 9175 23420
rect 9111 23360 9175 23364
rect 9191 23420 9255 23424
rect 9191 23364 9195 23420
rect 9195 23364 9251 23420
rect 9251 23364 9255 23420
rect 9191 23360 9255 23364
rect 9271 23420 9335 23424
rect 9271 23364 9275 23420
rect 9275 23364 9331 23420
rect 9331 23364 9335 23420
rect 9271 23360 9335 23364
rect 9351 23420 9415 23424
rect 9351 23364 9355 23420
rect 9355 23364 9411 23420
rect 9411 23364 9415 23420
rect 9351 23360 9415 23364
rect 4215 22876 4279 22880
rect 4215 22820 4219 22876
rect 4219 22820 4275 22876
rect 4275 22820 4279 22876
rect 4215 22816 4279 22820
rect 4295 22876 4359 22880
rect 4295 22820 4299 22876
rect 4299 22820 4355 22876
rect 4355 22820 4359 22876
rect 4295 22816 4359 22820
rect 4375 22876 4439 22880
rect 4375 22820 4379 22876
rect 4379 22820 4435 22876
rect 4435 22820 4439 22876
rect 4375 22816 4439 22820
rect 4455 22876 4519 22880
rect 4455 22820 4459 22876
rect 4459 22820 4515 22876
rect 4515 22820 4519 22876
rect 4455 22816 4519 22820
rect 7479 22876 7543 22880
rect 7479 22820 7483 22876
rect 7483 22820 7539 22876
rect 7539 22820 7543 22876
rect 7479 22816 7543 22820
rect 7559 22876 7623 22880
rect 7559 22820 7563 22876
rect 7563 22820 7619 22876
rect 7619 22820 7623 22876
rect 7559 22816 7623 22820
rect 7639 22876 7703 22880
rect 7639 22820 7643 22876
rect 7643 22820 7699 22876
rect 7699 22820 7703 22876
rect 7639 22816 7703 22820
rect 7719 22876 7783 22880
rect 7719 22820 7723 22876
rect 7723 22820 7779 22876
rect 7779 22820 7783 22876
rect 7719 22816 7783 22820
rect 2584 22332 2648 22336
rect 2584 22276 2588 22332
rect 2588 22276 2644 22332
rect 2644 22276 2648 22332
rect 2584 22272 2648 22276
rect 2664 22332 2728 22336
rect 2664 22276 2668 22332
rect 2668 22276 2724 22332
rect 2724 22276 2728 22332
rect 2664 22272 2728 22276
rect 2744 22332 2808 22336
rect 2744 22276 2748 22332
rect 2748 22276 2804 22332
rect 2804 22276 2808 22332
rect 2744 22272 2808 22276
rect 2824 22332 2888 22336
rect 2824 22276 2828 22332
rect 2828 22276 2884 22332
rect 2884 22276 2888 22332
rect 2824 22272 2888 22276
rect 5847 22332 5911 22336
rect 5847 22276 5851 22332
rect 5851 22276 5907 22332
rect 5907 22276 5911 22332
rect 5847 22272 5911 22276
rect 5927 22332 5991 22336
rect 5927 22276 5931 22332
rect 5931 22276 5987 22332
rect 5987 22276 5991 22332
rect 5927 22272 5991 22276
rect 6007 22332 6071 22336
rect 6007 22276 6011 22332
rect 6011 22276 6067 22332
rect 6067 22276 6071 22332
rect 6007 22272 6071 22276
rect 6087 22332 6151 22336
rect 6087 22276 6091 22332
rect 6091 22276 6147 22332
rect 6147 22276 6151 22332
rect 6087 22272 6151 22276
rect 9111 22332 9175 22336
rect 9111 22276 9115 22332
rect 9115 22276 9171 22332
rect 9171 22276 9175 22332
rect 9111 22272 9175 22276
rect 9191 22332 9255 22336
rect 9191 22276 9195 22332
rect 9195 22276 9251 22332
rect 9251 22276 9255 22332
rect 9191 22272 9255 22276
rect 9271 22332 9335 22336
rect 9271 22276 9275 22332
rect 9275 22276 9331 22332
rect 9331 22276 9335 22332
rect 9271 22272 9335 22276
rect 9351 22332 9415 22336
rect 9351 22276 9355 22332
rect 9355 22276 9411 22332
rect 9411 22276 9415 22332
rect 9351 22272 9415 22276
rect 4215 21788 4279 21792
rect 4215 21732 4219 21788
rect 4219 21732 4275 21788
rect 4275 21732 4279 21788
rect 4215 21728 4279 21732
rect 4295 21788 4359 21792
rect 4295 21732 4299 21788
rect 4299 21732 4355 21788
rect 4355 21732 4359 21788
rect 4295 21728 4359 21732
rect 4375 21788 4439 21792
rect 4375 21732 4379 21788
rect 4379 21732 4435 21788
rect 4435 21732 4439 21788
rect 4375 21728 4439 21732
rect 4455 21788 4519 21792
rect 4455 21732 4459 21788
rect 4459 21732 4515 21788
rect 4515 21732 4519 21788
rect 4455 21728 4519 21732
rect 7479 21788 7543 21792
rect 7479 21732 7483 21788
rect 7483 21732 7539 21788
rect 7539 21732 7543 21788
rect 7479 21728 7543 21732
rect 7559 21788 7623 21792
rect 7559 21732 7563 21788
rect 7563 21732 7619 21788
rect 7619 21732 7623 21788
rect 7559 21728 7623 21732
rect 7639 21788 7703 21792
rect 7639 21732 7643 21788
rect 7643 21732 7699 21788
rect 7699 21732 7703 21788
rect 7639 21728 7703 21732
rect 7719 21788 7783 21792
rect 7719 21732 7723 21788
rect 7723 21732 7779 21788
rect 7779 21732 7783 21788
rect 7719 21728 7783 21732
rect 2584 21244 2648 21248
rect 2584 21188 2588 21244
rect 2588 21188 2644 21244
rect 2644 21188 2648 21244
rect 2584 21184 2648 21188
rect 2664 21244 2728 21248
rect 2664 21188 2668 21244
rect 2668 21188 2724 21244
rect 2724 21188 2728 21244
rect 2664 21184 2728 21188
rect 2744 21244 2808 21248
rect 2744 21188 2748 21244
rect 2748 21188 2804 21244
rect 2804 21188 2808 21244
rect 2744 21184 2808 21188
rect 2824 21244 2888 21248
rect 2824 21188 2828 21244
rect 2828 21188 2884 21244
rect 2884 21188 2888 21244
rect 2824 21184 2888 21188
rect 5847 21244 5911 21248
rect 5847 21188 5851 21244
rect 5851 21188 5907 21244
rect 5907 21188 5911 21244
rect 5847 21184 5911 21188
rect 5927 21244 5991 21248
rect 5927 21188 5931 21244
rect 5931 21188 5987 21244
rect 5987 21188 5991 21244
rect 5927 21184 5991 21188
rect 6007 21244 6071 21248
rect 6007 21188 6011 21244
rect 6011 21188 6067 21244
rect 6067 21188 6071 21244
rect 6007 21184 6071 21188
rect 6087 21244 6151 21248
rect 6087 21188 6091 21244
rect 6091 21188 6147 21244
rect 6147 21188 6151 21244
rect 6087 21184 6151 21188
rect 9111 21244 9175 21248
rect 9111 21188 9115 21244
rect 9115 21188 9171 21244
rect 9171 21188 9175 21244
rect 9111 21184 9175 21188
rect 9191 21244 9255 21248
rect 9191 21188 9195 21244
rect 9195 21188 9251 21244
rect 9251 21188 9255 21244
rect 9191 21184 9255 21188
rect 9271 21244 9335 21248
rect 9271 21188 9275 21244
rect 9275 21188 9331 21244
rect 9331 21188 9335 21244
rect 9271 21184 9335 21188
rect 9351 21244 9415 21248
rect 9351 21188 9355 21244
rect 9355 21188 9411 21244
rect 9411 21188 9415 21244
rect 9351 21184 9415 21188
rect 4215 20700 4279 20704
rect 4215 20644 4219 20700
rect 4219 20644 4275 20700
rect 4275 20644 4279 20700
rect 4215 20640 4279 20644
rect 4295 20700 4359 20704
rect 4295 20644 4299 20700
rect 4299 20644 4355 20700
rect 4355 20644 4359 20700
rect 4295 20640 4359 20644
rect 4375 20700 4439 20704
rect 4375 20644 4379 20700
rect 4379 20644 4435 20700
rect 4435 20644 4439 20700
rect 4375 20640 4439 20644
rect 4455 20700 4519 20704
rect 4455 20644 4459 20700
rect 4459 20644 4515 20700
rect 4515 20644 4519 20700
rect 4455 20640 4519 20644
rect 7479 20700 7543 20704
rect 7479 20644 7483 20700
rect 7483 20644 7539 20700
rect 7539 20644 7543 20700
rect 7479 20640 7543 20644
rect 7559 20700 7623 20704
rect 7559 20644 7563 20700
rect 7563 20644 7619 20700
rect 7619 20644 7623 20700
rect 7559 20640 7623 20644
rect 7639 20700 7703 20704
rect 7639 20644 7643 20700
rect 7643 20644 7699 20700
rect 7699 20644 7703 20700
rect 7639 20640 7703 20644
rect 7719 20700 7783 20704
rect 7719 20644 7723 20700
rect 7723 20644 7779 20700
rect 7779 20644 7783 20700
rect 7719 20640 7783 20644
rect 2584 20156 2648 20160
rect 2584 20100 2588 20156
rect 2588 20100 2644 20156
rect 2644 20100 2648 20156
rect 2584 20096 2648 20100
rect 2664 20156 2728 20160
rect 2664 20100 2668 20156
rect 2668 20100 2724 20156
rect 2724 20100 2728 20156
rect 2664 20096 2728 20100
rect 2744 20156 2808 20160
rect 2744 20100 2748 20156
rect 2748 20100 2804 20156
rect 2804 20100 2808 20156
rect 2744 20096 2808 20100
rect 2824 20156 2888 20160
rect 2824 20100 2828 20156
rect 2828 20100 2884 20156
rect 2884 20100 2888 20156
rect 2824 20096 2888 20100
rect 5847 20156 5911 20160
rect 5847 20100 5851 20156
rect 5851 20100 5907 20156
rect 5907 20100 5911 20156
rect 5847 20096 5911 20100
rect 5927 20156 5991 20160
rect 5927 20100 5931 20156
rect 5931 20100 5987 20156
rect 5987 20100 5991 20156
rect 5927 20096 5991 20100
rect 6007 20156 6071 20160
rect 6007 20100 6011 20156
rect 6011 20100 6067 20156
rect 6067 20100 6071 20156
rect 6007 20096 6071 20100
rect 6087 20156 6151 20160
rect 6087 20100 6091 20156
rect 6091 20100 6147 20156
rect 6147 20100 6151 20156
rect 6087 20096 6151 20100
rect 9111 20156 9175 20160
rect 9111 20100 9115 20156
rect 9115 20100 9171 20156
rect 9171 20100 9175 20156
rect 9111 20096 9175 20100
rect 9191 20156 9255 20160
rect 9191 20100 9195 20156
rect 9195 20100 9251 20156
rect 9251 20100 9255 20156
rect 9191 20096 9255 20100
rect 9271 20156 9335 20160
rect 9271 20100 9275 20156
rect 9275 20100 9331 20156
rect 9331 20100 9335 20156
rect 9271 20096 9335 20100
rect 9351 20156 9415 20160
rect 9351 20100 9355 20156
rect 9355 20100 9411 20156
rect 9411 20100 9415 20156
rect 9351 20096 9415 20100
rect 4215 19612 4279 19616
rect 4215 19556 4219 19612
rect 4219 19556 4275 19612
rect 4275 19556 4279 19612
rect 4215 19552 4279 19556
rect 4295 19612 4359 19616
rect 4295 19556 4299 19612
rect 4299 19556 4355 19612
rect 4355 19556 4359 19612
rect 4295 19552 4359 19556
rect 4375 19612 4439 19616
rect 4375 19556 4379 19612
rect 4379 19556 4435 19612
rect 4435 19556 4439 19612
rect 4375 19552 4439 19556
rect 4455 19612 4519 19616
rect 4455 19556 4459 19612
rect 4459 19556 4515 19612
rect 4515 19556 4519 19612
rect 4455 19552 4519 19556
rect 7479 19612 7543 19616
rect 7479 19556 7483 19612
rect 7483 19556 7539 19612
rect 7539 19556 7543 19612
rect 7479 19552 7543 19556
rect 7559 19612 7623 19616
rect 7559 19556 7563 19612
rect 7563 19556 7619 19612
rect 7619 19556 7623 19612
rect 7559 19552 7623 19556
rect 7639 19612 7703 19616
rect 7639 19556 7643 19612
rect 7643 19556 7699 19612
rect 7699 19556 7703 19612
rect 7639 19552 7703 19556
rect 7719 19612 7783 19616
rect 7719 19556 7723 19612
rect 7723 19556 7779 19612
rect 7779 19556 7783 19612
rect 7719 19552 7783 19556
rect 2584 19068 2648 19072
rect 2584 19012 2588 19068
rect 2588 19012 2644 19068
rect 2644 19012 2648 19068
rect 2584 19008 2648 19012
rect 2664 19068 2728 19072
rect 2664 19012 2668 19068
rect 2668 19012 2724 19068
rect 2724 19012 2728 19068
rect 2664 19008 2728 19012
rect 2744 19068 2808 19072
rect 2744 19012 2748 19068
rect 2748 19012 2804 19068
rect 2804 19012 2808 19068
rect 2744 19008 2808 19012
rect 2824 19068 2888 19072
rect 2824 19012 2828 19068
rect 2828 19012 2884 19068
rect 2884 19012 2888 19068
rect 2824 19008 2888 19012
rect 5847 19068 5911 19072
rect 5847 19012 5851 19068
rect 5851 19012 5907 19068
rect 5907 19012 5911 19068
rect 5847 19008 5911 19012
rect 5927 19068 5991 19072
rect 5927 19012 5931 19068
rect 5931 19012 5987 19068
rect 5987 19012 5991 19068
rect 5927 19008 5991 19012
rect 6007 19068 6071 19072
rect 6007 19012 6011 19068
rect 6011 19012 6067 19068
rect 6067 19012 6071 19068
rect 6007 19008 6071 19012
rect 6087 19068 6151 19072
rect 6087 19012 6091 19068
rect 6091 19012 6147 19068
rect 6147 19012 6151 19068
rect 6087 19008 6151 19012
rect 9111 19068 9175 19072
rect 9111 19012 9115 19068
rect 9115 19012 9171 19068
rect 9171 19012 9175 19068
rect 9111 19008 9175 19012
rect 9191 19068 9255 19072
rect 9191 19012 9195 19068
rect 9195 19012 9251 19068
rect 9251 19012 9255 19068
rect 9191 19008 9255 19012
rect 9271 19068 9335 19072
rect 9271 19012 9275 19068
rect 9275 19012 9331 19068
rect 9331 19012 9335 19068
rect 9271 19008 9335 19012
rect 9351 19068 9415 19072
rect 9351 19012 9355 19068
rect 9355 19012 9411 19068
rect 9411 19012 9415 19068
rect 9351 19008 9415 19012
rect 4215 18524 4279 18528
rect 4215 18468 4219 18524
rect 4219 18468 4275 18524
rect 4275 18468 4279 18524
rect 4215 18464 4279 18468
rect 4295 18524 4359 18528
rect 4295 18468 4299 18524
rect 4299 18468 4355 18524
rect 4355 18468 4359 18524
rect 4295 18464 4359 18468
rect 4375 18524 4439 18528
rect 4375 18468 4379 18524
rect 4379 18468 4435 18524
rect 4435 18468 4439 18524
rect 4375 18464 4439 18468
rect 4455 18524 4519 18528
rect 4455 18468 4459 18524
rect 4459 18468 4515 18524
rect 4515 18468 4519 18524
rect 4455 18464 4519 18468
rect 7479 18524 7543 18528
rect 7479 18468 7483 18524
rect 7483 18468 7539 18524
rect 7539 18468 7543 18524
rect 7479 18464 7543 18468
rect 7559 18524 7623 18528
rect 7559 18468 7563 18524
rect 7563 18468 7619 18524
rect 7619 18468 7623 18524
rect 7559 18464 7623 18468
rect 7639 18524 7703 18528
rect 7639 18468 7643 18524
rect 7643 18468 7699 18524
rect 7699 18468 7703 18524
rect 7639 18464 7703 18468
rect 7719 18524 7783 18528
rect 7719 18468 7723 18524
rect 7723 18468 7779 18524
rect 7779 18468 7783 18524
rect 7719 18464 7783 18468
rect 2584 17980 2648 17984
rect 2584 17924 2588 17980
rect 2588 17924 2644 17980
rect 2644 17924 2648 17980
rect 2584 17920 2648 17924
rect 2664 17980 2728 17984
rect 2664 17924 2668 17980
rect 2668 17924 2724 17980
rect 2724 17924 2728 17980
rect 2664 17920 2728 17924
rect 2744 17980 2808 17984
rect 2744 17924 2748 17980
rect 2748 17924 2804 17980
rect 2804 17924 2808 17980
rect 2744 17920 2808 17924
rect 2824 17980 2888 17984
rect 2824 17924 2828 17980
rect 2828 17924 2884 17980
rect 2884 17924 2888 17980
rect 2824 17920 2888 17924
rect 5847 17980 5911 17984
rect 5847 17924 5851 17980
rect 5851 17924 5907 17980
rect 5907 17924 5911 17980
rect 5847 17920 5911 17924
rect 5927 17980 5991 17984
rect 5927 17924 5931 17980
rect 5931 17924 5987 17980
rect 5987 17924 5991 17980
rect 5927 17920 5991 17924
rect 6007 17980 6071 17984
rect 6007 17924 6011 17980
rect 6011 17924 6067 17980
rect 6067 17924 6071 17980
rect 6007 17920 6071 17924
rect 6087 17980 6151 17984
rect 6087 17924 6091 17980
rect 6091 17924 6147 17980
rect 6147 17924 6151 17980
rect 6087 17920 6151 17924
rect 9111 17980 9175 17984
rect 9111 17924 9115 17980
rect 9115 17924 9171 17980
rect 9171 17924 9175 17980
rect 9111 17920 9175 17924
rect 9191 17980 9255 17984
rect 9191 17924 9195 17980
rect 9195 17924 9251 17980
rect 9251 17924 9255 17980
rect 9191 17920 9255 17924
rect 9271 17980 9335 17984
rect 9271 17924 9275 17980
rect 9275 17924 9331 17980
rect 9331 17924 9335 17980
rect 9271 17920 9335 17924
rect 9351 17980 9415 17984
rect 9351 17924 9355 17980
rect 9355 17924 9411 17980
rect 9411 17924 9415 17980
rect 9351 17920 9415 17924
rect 4215 17436 4279 17440
rect 4215 17380 4219 17436
rect 4219 17380 4275 17436
rect 4275 17380 4279 17436
rect 4215 17376 4279 17380
rect 4295 17436 4359 17440
rect 4295 17380 4299 17436
rect 4299 17380 4355 17436
rect 4355 17380 4359 17436
rect 4295 17376 4359 17380
rect 4375 17436 4439 17440
rect 4375 17380 4379 17436
rect 4379 17380 4435 17436
rect 4435 17380 4439 17436
rect 4375 17376 4439 17380
rect 4455 17436 4519 17440
rect 4455 17380 4459 17436
rect 4459 17380 4515 17436
rect 4515 17380 4519 17436
rect 4455 17376 4519 17380
rect 7479 17436 7543 17440
rect 7479 17380 7483 17436
rect 7483 17380 7539 17436
rect 7539 17380 7543 17436
rect 7479 17376 7543 17380
rect 7559 17436 7623 17440
rect 7559 17380 7563 17436
rect 7563 17380 7619 17436
rect 7619 17380 7623 17436
rect 7559 17376 7623 17380
rect 7639 17436 7703 17440
rect 7639 17380 7643 17436
rect 7643 17380 7699 17436
rect 7699 17380 7703 17436
rect 7639 17376 7703 17380
rect 7719 17436 7783 17440
rect 7719 17380 7723 17436
rect 7723 17380 7779 17436
rect 7779 17380 7783 17436
rect 7719 17376 7783 17380
rect 2584 16892 2648 16896
rect 2584 16836 2588 16892
rect 2588 16836 2644 16892
rect 2644 16836 2648 16892
rect 2584 16832 2648 16836
rect 2664 16892 2728 16896
rect 2664 16836 2668 16892
rect 2668 16836 2724 16892
rect 2724 16836 2728 16892
rect 2664 16832 2728 16836
rect 2744 16892 2808 16896
rect 2744 16836 2748 16892
rect 2748 16836 2804 16892
rect 2804 16836 2808 16892
rect 2744 16832 2808 16836
rect 2824 16892 2888 16896
rect 2824 16836 2828 16892
rect 2828 16836 2884 16892
rect 2884 16836 2888 16892
rect 2824 16832 2888 16836
rect 5847 16892 5911 16896
rect 5847 16836 5851 16892
rect 5851 16836 5907 16892
rect 5907 16836 5911 16892
rect 5847 16832 5911 16836
rect 5927 16892 5991 16896
rect 5927 16836 5931 16892
rect 5931 16836 5987 16892
rect 5987 16836 5991 16892
rect 5927 16832 5991 16836
rect 6007 16892 6071 16896
rect 6007 16836 6011 16892
rect 6011 16836 6067 16892
rect 6067 16836 6071 16892
rect 6007 16832 6071 16836
rect 6087 16892 6151 16896
rect 6087 16836 6091 16892
rect 6091 16836 6147 16892
rect 6147 16836 6151 16892
rect 6087 16832 6151 16836
rect 9111 16892 9175 16896
rect 9111 16836 9115 16892
rect 9115 16836 9171 16892
rect 9171 16836 9175 16892
rect 9111 16832 9175 16836
rect 9191 16892 9255 16896
rect 9191 16836 9195 16892
rect 9195 16836 9251 16892
rect 9251 16836 9255 16892
rect 9191 16832 9255 16836
rect 9271 16892 9335 16896
rect 9271 16836 9275 16892
rect 9275 16836 9331 16892
rect 9331 16836 9335 16892
rect 9271 16832 9335 16836
rect 9351 16892 9415 16896
rect 9351 16836 9355 16892
rect 9355 16836 9411 16892
rect 9411 16836 9415 16892
rect 9351 16832 9415 16836
rect 4215 16348 4279 16352
rect 4215 16292 4219 16348
rect 4219 16292 4275 16348
rect 4275 16292 4279 16348
rect 4215 16288 4279 16292
rect 4295 16348 4359 16352
rect 4295 16292 4299 16348
rect 4299 16292 4355 16348
rect 4355 16292 4359 16348
rect 4295 16288 4359 16292
rect 4375 16348 4439 16352
rect 4375 16292 4379 16348
rect 4379 16292 4435 16348
rect 4435 16292 4439 16348
rect 4375 16288 4439 16292
rect 4455 16348 4519 16352
rect 4455 16292 4459 16348
rect 4459 16292 4515 16348
rect 4515 16292 4519 16348
rect 4455 16288 4519 16292
rect 7479 16348 7543 16352
rect 7479 16292 7483 16348
rect 7483 16292 7539 16348
rect 7539 16292 7543 16348
rect 7479 16288 7543 16292
rect 7559 16348 7623 16352
rect 7559 16292 7563 16348
rect 7563 16292 7619 16348
rect 7619 16292 7623 16348
rect 7559 16288 7623 16292
rect 7639 16348 7703 16352
rect 7639 16292 7643 16348
rect 7643 16292 7699 16348
rect 7699 16292 7703 16348
rect 7639 16288 7703 16292
rect 7719 16348 7783 16352
rect 7719 16292 7723 16348
rect 7723 16292 7779 16348
rect 7779 16292 7783 16348
rect 7719 16288 7783 16292
rect 2584 15804 2648 15808
rect 2584 15748 2588 15804
rect 2588 15748 2644 15804
rect 2644 15748 2648 15804
rect 2584 15744 2648 15748
rect 2664 15804 2728 15808
rect 2664 15748 2668 15804
rect 2668 15748 2724 15804
rect 2724 15748 2728 15804
rect 2664 15744 2728 15748
rect 2744 15804 2808 15808
rect 2744 15748 2748 15804
rect 2748 15748 2804 15804
rect 2804 15748 2808 15804
rect 2744 15744 2808 15748
rect 2824 15804 2888 15808
rect 2824 15748 2828 15804
rect 2828 15748 2884 15804
rect 2884 15748 2888 15804
rect 2824 15744 2888 15748
rect 5847 15804 5911 15808
rect 5847 15748 5851 15804
rect 5851 15748 5907 15804
rect 5907 15748 5911 15804
rect 5847 15744 5911 15748
rect 5927 15804 5991 15808
rect 5927 15748 5931 15804
rect 5931 15748 5987 15804
rect 5987 15748 5991 15804
rect 5927 15744 5991 15748
rect 6007 15804 6071 15808
rect 6007 15748 6011 15804
rect 6011 15748 6067 15804
rect 6067 15748 6071 15804
rect 6007 15744 6071 15748
rect 6087 15804 6151 15808
rect 6087 15748 6091 15804
rect 6091 15748 6147 15804
rect 6147 15748 6151 15804
rect 6087 15744 6151 15748
rect 9111 15804 9175 15808
rect 9111 15748 9115 15804
rect 9115 15748 9171 15804
rect 9171 15748 9175 15804
rect 9111 15744 9175 15748
rect 9191 15804 9255 15808
rect 9191 15748 9195 15804
rect 9195 15748 9251 15804
rect 9251 15748 9255 15804
rect 9191 15744 9255 15748
rect 9271 15804 9335 15808
rect 9271 15748 9275 15804
rect 9275 15748 9331 15804
rect 9331 15748 9335 15804
rect 9271 15744 9335 15748
rect 9351 15804 9415 15808
rect 9351 15748 9355 15804
rect 9355 15748 9411 15804
rect 9411 15748 9415 15804
rect 9351 15744 9415 15748
rect 4215 15260 4279 15264
rect 4215 15204 4219 15260
rect 4219 15204 4275 15260
rect 4275 15204 4279 15260
rect 4215 15200 4279 15204
rect 4295 15260 4359 15264
rect 4295 15204 4299 15260
rect 4299 15204 4355 15260
rect 4355 15204 4359 15260
rect 4295 15200 4359 15204
rect 4375 15260 4439 15264
rect 4375 15204 4379 15260
rect 4379 15204 4435 15260
rect 4435 15204 4439 15260
rect 4375 15200 4439 15204
rect 4455 15260 4519 15264
rect 4455 15204 4459 15260
rect 4459 15204 4515 15260
rect 4515 15204 4519 15260
rect 4455 15200 4519 15204
rect 7479 15260 7543 15264
rect 7479 15204 7483 15260
rect 7483 15204 7539 15260
rect 7539 15204 7543 15260
rect 7479 15200 7543 15204
rect 7559 15260 7623 15264
rect 7559 15204 7563 15260
rect 7563 15204 7619 15260
rect 7619 15204 7623 15260
rect 7559 15200 7623 15204
rect 7639 15260 7703 15264
rect 7639 15204 7643 15260
rect 7643 15204 7699 15260
rect 7699 15204 7703 15260
rect 7639 15200 7703 15204
rect 7719 15260 7783 15264
rect 7719 15204 7723 15260
rect 7723 15204 7779 15260
rect 7779 15204 7783 15260
rect 7719 15200 7783 15204
rect 2584 14716 2648 14720
rect 2584 14660 2588 14716
rect 2588 14660 2644 14716
rect 2644 14660 2648 14716
rect 2584 14656 2648 14660
rect 2664 14716 2728 14720
rect 2664 14660 2668 14716
rect 2668 14660 2724 14716
rect 2724 14660 2728 14716
rect 2664 14656 2728 14660
rect 2744 14716 2808 14720
rect 2744 14660 2748 14716
rect 2748 14660 2804 14716
rect 2804 14660 2808 14716
rect 2744 14656 2808 14660
rect 2824 14716 2888 14720
rect 2824 14660 2828 14716
rect 2828 14660 2884 14716
rect 2884 14660 2888 14716
rect 2824 14656 2888 14660
rect 5847 14716 5911 14720
rect 5847 14660 5851 14716
rect 5851 14660 5907 14716
rect 5907 14660 5911 14716
rect 5847 14656 5911 14660
rect 5927 14716 5991 14720
rect 5927 14660 5931 14716
rect 5931 14660 5987 14716
rect 5987 14660 5991 14716
rect 5927 14656 5991 14660
rect 6007 14716 6071 14720
rect 6007 14660 6011 14716
rect 6011 14660 6067 14716
rect 6067 14660 6071 14716
rect 6007 14656 6071 14660
rect 6087 14716 6151 14720
rect 6087 14660 6091 14716
rect 6091 14660 6147 14716
rect 6147 14660 6151 14716
rect 6087 14656 6151 14660
rect 9111 14716 9175 14720
rect 9111 14660 9115 14716
rect 9115 14660 9171 14716
rect 9171 14660 9175 14716
rect 9111 14656 9175 14660
rect 9191 14716 9255 14720
rect 9191 14660 9195 14716
rect 9195 14660 9251 14716
rect 9251 14660 9255 14716
rect 9191 14656 9255 14660
rect 9271 14716 9335 14720
rect 9271 14660 9275 14716
rect 9275 14660 9331 14716
rect 9331 14660 9335 14716
rect 9271 14656 9335 14660
rect 9351 14716 9415 14720
rect 9351 14660 9355 14716
rect 9355 14660 9411 14716
rect 9411 14660 9415 14716
rect 9351 14656 9415 14660
rect 4215 14172 4279 14176
rect 4215 14116 4219 14172
rect 4219 14116 4275 14172
rect 4275 14116 4279 14172
rect 4215 14112 4279 14116
rect 4295 14172 4359 14176
rect 4295 14116 4299 14172
rect 4299 14116 4355 14172
rect 4355 14116 4359 14172
rect 4295 14112 4359 14116
rect 4375 14172 4439 14176
rect 4375 14116 4379 14172
rect 4379 14116 4435 14172
rect 4435 14116 4439 14172
rect 4375 14112 4439 14116
rect 4455 14172 4519 14176
rect 4455 14116 4459 14172
rect 4459 14116 4515 14172
rect 4515 14116 4519 14172
rect 4455 14112 4519 14116
rect 7479 14172 7543 14176
rect 7479 14116 7483 14172
rect 7483 14116 7539 14172
rect 7539 14116 7543 14172
rect 7479 14112 7543 14116
rect 7559 14172 7623 14176
rect 7559 14116 7563 14172
rect 7563 14116 7619 14172
rect 7619 14116 7623 14172
rect 7559 14112 7623 14116
rect 7639 14172 7703 14176
rect 7639 14116 7643 14172
rect 7643 14116 7699 14172
rect 7699 14116 7703 14172
rect 7639 14112 7703 14116
rect 7719 14172 7783 14176
rect 7719 14116 7723 14172
rect 7723 14116 7779 14172
rect 7779 14116 7783 14172
rect 7719 14112 7783 14116
rect 2584 13628 2648 13632
rect 2584 13572 2588 13628
rect 2588 13572 2644 13628
rect 2644 13572 2648 13628
rect 2584 13568 2648 13572
rect 2664 13628 2728 13632
rect 2664 13572 2668 13628
rect 2668 13572 2724 13628
rect 2724 13572 2728 13628
rect 2664 13568 2728 13572
rect 2744 13628 2808 13632
rect 2744 13572 2748 13628
rect 2748 13572 2804 13628
rect 2804 13572 2808 13628
rect 2744 13568 2808 13572
rect 2824 13628 2888 13632
rect 2824 13572 2828 13628
rect 2828 13572 2884 13628
rect 2884 13572 2888 13628
rect 2824 13568 2888 13572
rect 5847 13628 5911 13632
rect 5847 13572 5851 13628
rect 5851 13572 5907 13628
rect 5907 13572 5911 13628
rect 5847 13568 5911 13572
rect 5927 13628 5991 13632
rect 5927 13572 5931 13628
rect 5931 13572 5987 13628
rect 5987 13572 5991 13628
rect 5927 13568 5991 13572
rect 6007 13628 6071 13632
rect 6007 13572 6011 13628
rect 6011 13572 6067 13628
rect 6067 13572 6071 13628
rect 6007 13568 6071 13572
rect 6087 13628 6151 13632
rect 6087 13572 6091 13628
rect 6091 13572 6147 13628
rect 6147 13572 6151 13628
rect 6087 13568 6151 13572
rect 9111 13628 9175 13632
rect 9111 13572 9115 13628
rect 9115 13572 9171 13628
rect 9171 13572 9175 13628
rect 9111 13568 9175 13572
rect 9191 13628 9255 13632
rect 9191 13572 9195 13628
rect 9195 13572 9251 13628
rect 9251 13572 9255 13628
rect 9191 13568 9255 13572
rect 9271 13628 9335 13632
rect 9271 13572 9275 13628
rect 9275 13572 9331 13628
rect 9331 13572 9335 13628
rect 9271 13568 9335 13572
rect 9351 13628 9415 13632
rect 9351 13572 9355 13628
rect 9355 13572 9411 13628
rect 9411 13572 9415 13628
rect 9351 13568 9415 13572
rect 4215 13084 4279 13088
rect 4215 13028 4219 13084
rect 4219 13028 4275 13084
rect 4275 13028 4279 13084
rect 4215 13024 4279 13028
rect 4295 13084 4359 13088
rect 4295 13028 4299 13084
rect 4299 13028 4355 13084
rect 4355 13028 4359 13084
rect 4295 13024 4359 13028
rect 4375 13084 4439 13088
rect 4375 13028 4379 13084
rect 4379 13028 4435 13084
rect 4435 13028 4439 13084
rect 4375 13024 4439 13028
rect 4455 13084 4519 13088
rect 4455 13028 4459 13084
rect 4459 13028 4515 13084
rect 4515 13028 4519 13084
rect 4455 13024 4519 13028
rect 7479 13084 7543 13088
rect 7479 13028 7483 13084
rect 7483 13028 7539 13084
rect 7539 13028 7543 13084
rect 7479 13024 7543 13028
rect 7559 13084 7623 13088
rect 7559 13028 7563 13084
rect 7563 13028 7619 13084
rect 7619 13028 7623 13084
rect 7559 13024 7623 13028
rect 7639 13084 7703 13088
rect 7639 13028 7643 13084
rect 7643 13028 7699 13084
rect 7699 13028 7703 13084
rect 7639 13024 7703 13028
rect 7719 13084 7783 13088
rect 7719 13028 7723 13084
rect 7723 13028 7779 13084
rect 7779 13028 7783 13084
rect 7719 13024 7783 13028
rect 2584 12540 2648 12544
rect 2584 12484 2588 12540
rect 2588 12484 2644 12540
rect 2644 12484 2648 12540
rect 2584 12480 2648 12484
rect 2664 12540 2728 12544
rect 2664 12484 2668 12540
rect 2668 12484 2724 12540
rect 2724 12484 2728 12540
rect 2664 12480 2728 12484
rect 2744 12540 2808 12544
rect 2744 12484 2748 12540
rect 2748 12484 2804 12540
rect 2804 12484 2808 12540
rect 2744 12480 2808 12484
rect 2824 12540 2888 12544
rect 2824 12484 2828 12540
rect 2828 12484 2884 12540
rect 2884 12484 2888 12540
rect 2824 12480 2888 12484
rect 5847 12540 5911 12544
rect 5847 12484 5851 12540
rect 5851 12484 5907 12540
rect 5907 12484 5911 12540
rect 5847 12480 5911 12484
rect 5927 12540 5991 12544
rect 5927 12484 5931 12540
rect 5931 12484 5987 12540
rect 5987 12484 5991 12540
rect 5927 12480 5991 12484
rect 6007 12540 6071 12544
rect 6007 12484 6011 12540
rect 6011 12484 6067 12540
rect 6067 12484 6071 12540
rect 6007 12480 6071 12484
rect 6087 12540 6151 12544
rect 6087 12484 6091 12540
rect 6091 12484 6147 12540
rect 6147 12484 6151 12540
rect 6087 12480 6151 12484
rect 9111 12540 9175 12544
rect 9111 12484 9115 12540
rect 9115 12484 9171 12540
rect 9171 12484 9175 12540
rect 9111 12480 9175 12484
rect 9191 12540 9255 12544
rect 9191 12484 9195 12540
rect 9195 12484 9251 12540
rect 9251 12484 9255 12540
rect 9191 12480 9255 12484
rect 9271 12540 9335 12544
rect 9271 12484 9275 12540
rect 9275 12484 9331 12540
rect 9331 12484 9335 12540
rect 9271 12480 9335 12484
rect 9351 12540 9415 12544
rect 9351 12484 9355 12540
rect 9355 12484 9411 12540
rect 9411 12484 9415 12540
rect 9351 12480 9415 12484
rect 4215 11996 4279 12000
rect 4215 11940 4219 11996
rect 4219 11940 4275 11996
rect 4275 11940 4279 11996
rect 4215 11936 4279 11940
rect 4295 11996 4359 12000
rect 4295 11940 4299 11996
rect 4299 11940 4355 11996
rect 4355 11940 4359 11996
rect 4295 11936 4359 11940
rect 4375 11996 4439 12000
rect 4375 11940 4379 11996
rect 4379 11940 4435 11996
rect 4435 11940 4439 11996
rect 4375 11936 4439 11940
rect 4455 11996 4519 12000
rect 4455 11940 4459 11996
rect 4459 11940 4515 11996
rect 4515 11940 4519 11996
rect 4455 11936 4519 11940
rect 7479 11996 7543 12000
rect 7479 11940 7483 11996
rect 7483 11940 7539 11996
rect 7539 11940 7543 11996
rect 7479 11936 7543 11940
rect 7559 11996 7623 12000
rect 7559 11940 7563 11996
rect 7563 11940 7619 11996
rect 7619 11940 7623 11996
rect 7559 11936 7623 11940
rect 7639 11996 7703 12000
rect 7639 11940 7643 11996
rect 7643 11940 7699 11996
rect 7699 11940 7703 11996
rect 7639 11936 7703 11940
rect 7719 11996 7783 12000
rect 7719 11940 7723 11996
rect 7723 11940 7779 11996
rect 7779 11940 7783 11996
rect 7719 11936 7783 11940
rect 2584 11452 2648 11456
rect 2584 11396 2588 11452
rect 2588 11396 2644 11452
rect 2644 11396 2648 11452
rect 2584 11392 2648 11396
rect 2664 11452 2728 11456
rect 2664 11396 2668 11452
rect 2668 11396 2724 11452
rect 2724 11396 2728 11452
rect 2664 11392 2728 11396
rect 2744 11452 2808 11456
rect 2744 11396 2748 11452
rect 2748 11396 2804 11452
rect 2804 11396 2808 11452
rect 2744 11392 2808 11396
rect 2824 11452 2888 11456
rect 2824 11396 2828 11452
rect 2828 11396 2884 11452
rect 2884 11396 2888 11452
rect 2824 11392 2888 11396
rect 5847 11452 5911 11456
rect 5847 11396 5851 11452
rect 5851 11396 5907 11452
rect 5907 11396 5911 11452
rect 5847 11392 5911 11396
rect 5927 11452 5991 11456
rect 5927 11396 5931 11452
rect 5931 11396 5987 11452
rect 5987 11396 5991 11452
rect 5927 11392 5991 11396
rect 6007 11452 6071 11456
rect 6007 11396 6011 11452
rect 6011 11396 6067 11452
rect 6067 11396 6071 11452
rect 6007 11392 6071 11396
rect 6087 11452 6151 11456
rect 6087 11396 6091 11452
rect 6091 11396 6147 11452
rect 6147 11396 6151 11452
rect 6087 11392 6151 11396
rect 9111 11452 9175 11456
rect 9111 11396 9115 11452
rect 9115 11396 9171 11452
rect 9171 11396 9175 11452
rect 9111 11392 9175 11396
rect 9191 11452 9255 11456
rect 9191 11396 9195 11452
rect 9195 11396 9251 11452
rect 9251 11396 9255 11452
rect 9191 11392 9255 11396
rect 9271 11452 9335 11456
rect 9271 11396 9275 11452
rect 9275 11396 9331 11452
rect 9331 11396 9335 11452
rect 9271 11392 9335 11396
rect 9351 11452 9415 11456
rect 9351 11396 9355 11452
rect 9355 11396 9411 11452
rect 9411 11396 9415 11452
rect 9351 11392 9415 11396
rect 4215 10908 4279 10912
rect 4215 10852 4219 10908
rect 4219 10852 4275 10908
rect 4275 10852 4279 10908
rect 4215 10848 4279 10852
rect 4295 10908 4359 10912
rect 4295 10852 4299 10908
rect 4299 10852 4355 10908
rect 4355 10852 4359 10908
rect 4295 10848 4359 10852
rect 4375 10908 4439 10912
rect 4375 10852 4379 10908
rect 4379 10852 4435 10908
rect 4435 10852 4439 10908
rect 4375 10848 4439 10852
rect 4455 10908 4519 10912
rect 4455 10852 4459 10908
rect 4459 10852 4515 10908
rect 4515 10852 4519 10908
rect 4455 10848 4519 10852
rect 7479 10908 7543 10912
rect 7479 10852 7483 10908
rect 7483 10852 7539 10908
rect 7539 10852 7543 10908
rect 7479 10848 7543 10852
rect 7559 10908 7623 10912
rect 7559 10852 7563 10908
rect 7563 10852 7619 10908
rect 7619 10852 7623 10908
rect 7559 10848 7623 10852
rect 7639 10908 7703 10912
rect 7639 10852 7643 10908
rect 7643 10852 7699 10908
rect 7699 10852 7703 10908
rect 7639 10848 7703 10852
rect 7719 10908 7783 10912
rect 7719 10852 7723 10908
rect 7723 10852 7779 10908
rect 7779 10852 7783 10908
rect 7719 10848 7783 10852
rect 2584 10364 2648 10368
rect 2584 10308 2588 10364
rect 2588 10308 2644 10364
rect 2644 10308 2648 10364
rect 2584 10304 2648 10308
rect 2664 10364 2728 10368
rect 2664 10308 2668 10364
rect 2668 10308 2724 10364
rect 2724 10308 2728 10364
rect 2664 10304 2728 10308
rect 2744 10364 2808 10368
rect 2744 10308 2748 10364
rect 2748 10308 2804 10364
rect 2804 10308 2808 10364
rect 2744 10304 2808 10308
rect 2824 10364 2888 10368
rect 2824 10308 2828 10364
rect 2828 10308 2884 10364
rect 2884 10308 2888 10364
rect 2824 10304 2888 10308
rect 5847 10364 5911 10368
rect 5847 10308 5851 10364
rect 5851 10308 5907 10364
rect 5907 10308 5911 10364
rect 5847 10304 5911 10308
rect 5927 10364 5991 10368
rect 5927 10308 5931 10364
rect 5931 10308 5987 10364
rect 5987 10308 5991 10364
rect 5927 10304 5991 10308
rect 6007 10364 6071 10368
rect 6007 10308 6011 10364
rect 6011 10308 6067 10364
rect 6067 10308 6071 10364
rect 6007 10304 6071 10308
rect 6087 10364 6151 10368
rect 6087 10308 6091 10364
rect 6091 10308 6147 10364
rect 6147 10308 6151 10364
rect 6087 10304 6151 10308
rect 9111 10364 9175 10368
rect 9111 10308 9115 10364
rect 9115 10308 9171 10364
rect 9171 10308 9175 10364
rect 9111 10304 9175 10308
rect 9191 10364 9255 10368
rect 9191 10308 9195 10364
rect 9195 10308 9251 10364
rect 9251 10308 9255 10364
rect 9191 10304 9255 10308
rect 9271 10364 9335 10368
rect 9271 10308 9275 10364
rect 9275 10308 9331 10364
rect 9331 10308 9335 10364
rect 9271 10304 9335 10308
rect 9351 10364 9415 10368
rect 9351 10308 9355 10364
rect 9355 10308 9411 10364
rect 9411 10308 9415 10364
rect 9351 10304 9415 10308
rect 4215 9820 4279 9824
rect 4215 9764 4219 9820
rect 4219 9764 4275 9820
rect 4275 9764 4279 9820
rect 4215 9760 4279 9764
rect 4295 9820 4359 9824
rect 4295 9764 4299 9820
rect 4299 9764 4355 9820
rect 4355 9764 4359 9820
rect 4295 9760 4359 9764
rect 4375 9820 4439 9824
rect 4375 9764 4379 9820
rect 4379 9764 4435 9820
rect 4435 9764 4439 9820
rect 4375 9760 4439 9764
rect 4455 9820 4519 9824
rect 4455 9764 4459 9820
rect 4459 9764 4515 9820
rect 4515 9764 4519 9820
rect 4455 9760 4519 9764
rect 7479 9820 7543 9824
rect 7479 9764 7483 9820
rect 7483 9764 7539 9820
rect 7539 9764 7543 9820
rect 7479 9760 7543 9764
rect 7559 9820 7623 9824
rect 7559 9764 7563 9820
rect 7563 9764 7619 9820
rect 7619 9764 7623 9820
rect 7559 9760 7623 9764
rect 7639 9820 7703 9824
rect 7639 9764 7643 9820
rect 7643 9764 7699 9820
rect 7699 9764 7703 9820
rect 7639 9760 7703 9764
rect 7719 9820 7783 9824
rect 7719 9764 7723 9820
rect 7723 9764 7779 9820
rect 7779 9764 7783 9820
rect 7719 9760 7783 9764
rect 2584 9276 2648 9280
rect 2584 9220 2588 9276
rect 2588 9220 2644 9276
rect 2644 9220 2648 9276
rect 2584 9216 2648 9220
rect 2664 9276 2728 9280
rect 2664 9220 2668 9276
rect 2668 9220 2724 9276
rect 2724 9220 2728 9276
rect 2664 9216 2728 9220
rect 2744 9276 2808 9280
rect 2744 9220 2748 9276
rect 2748 9220 2804 9276
rect 2804 9220 2808 9276
rect 2744 9216 2808 9220
rect 2824 9276 2888 9280
rect 2824 9220 2828 9276
rect 2828 9220 2884 9276
rect 2884 9220 2888 9276
rect 2824 9216 2888 9220
rect 5847 9276 5911 9280
rect 5847 9220 5851 9276
rect 5851 9220 5907 9276
rect 5907 9220 5911 9276
rect 5847 9216 5911 9220
rect 5927 9276 5991 9280
rect 5927 9220 5931 9276
rect 5931 9220 5987 9276
rect 5987 9220 5991 9276
rect 5927 9216 5991 9220
rect 6007 9276 6071 9280
rect 6007 9220 6011 9276
rect 6011 9220 6067 9276
rect 6067 9220 6071 9276
rect 6007 9216 6071 9220
rect 6087 9276 6151 9280
rect 6087 9220 6091 9276
rect 6091 9220 6147 9276
rect 6147 9220 6151 9276
rect 6087 9216 6151 9220
rect 9111 9276 9175 9280
rect 9111 9220 9115 9276
rect 9115 9220 9171 9276
rect 9171 9220 9175 9276
rect 9111 9216 9175 9220
rect 9191 9276 9255 9280
rect 9191 9220 9195 9276
rect 9195 9220 9251 9276
rect 9251 9220 9255 9276
rect 9191 9216 9255 9220
rect 9271 9276 9335 9280
rect 9271 9220 9275 9276
rect 9275 9220 9331 9276
rect 9331 9220 9335 9276
rect 9271 9216 9335 9220
rect 9351 9276 9415 9280
rect 9351 9220 9355 9276
rect 9355 9220 9411 9276
rect 9411 9220 9415 9276
rect 9351 9216 9415 9220
rect 4215 8732 4279 8736
rect 4215 8676 4219 8732
rect 4219 8676 4275 8732
rect 4275 8676 4279 8732
rect 4215 8672 4279 8676
rect 4295 8732 4359 8736
rect 4295 8676 4299 8732
rect 4299 8676 4355 8732
rect 4355 8676 4359 8732
rect 4295 8672 4359 8676
rect 4375 8732 4439 8736
rect 4375 8676 4379 8732
rect 4379 8676 4435 8732
rect 4435 8676 4439 8732
rect 4375 8672 4439 8676
rect 4455 8732 4519 8736
rect 4455 8676 4459 8732
rect 4459 8676 4515 8732
rect 4515 8676 4519 8732
rect 4455 8672 4519 8676
rect 7479 8732 7543 8736
rect 7479 8676 7483 8732
rect 7483 8676 7539 8732
rect 7539 8676 7543 8732
rect 7479 8672 7543 8676
rect 7559 8732 7623 8736
rect 7559 8676 7563 8732
rect 7563 8676 7619 8732
rect 7619 8676 7623 8732
rect 7559 8672 7623 8676
rect 7639 8732 7703 8736
rect 7639 8676 7643 8732
rect 7643 8676 7699 8732
rect 7699 8676 7703 8732
rect 7639 8672 7703 8676
rect 7719 8732 7783 8736
rect 7719 8676 7723 8732
rect 7723 8676 7779 8732
rect 7779 8676 7783 8732
rect 7719 8672 7783 8676
rect 2584 8188 2648 8192
rect 2584 8132 2588 8188
rect 2588 8132 2644 8188
rect 2644 8132 2648 8188
rect 2584 8128 2648 8132
rect 2664 8188 2728 8192
rect 2664 8132 2668 8188
rect 2668 8132 2724 8188
rect 2724 8132 2728 8188
rect 2664 8128 2728 8132
rect 2744 8188 2808 8192
rect 2744 8132 2748 8188
rect 2748 8132 2804 8188
rect 2804 8132 2808 8188
rect 2744 8128 2808 8132
rect 2824 8188 2888 8192
rect 2824 8132 2828 8188
rect 2828 8132 2884 8188
rect 2884 8132 2888 8188
rect 2824 8128 2888 8132
rect 5847 8188 5911 8192
rect 5847 8132 5851 8188
rect 5851 8132 5907 8188
rect 5907 8132 5911 8188
rect 5847 8128 5911 8132
rect 5927 8188 5991 8192
rect 5927 8132 5931 8188
rect 5931 8132 5987 8188
rect 5987 8132 5991 8188
rect 5927 8128 5991 8132
rect 6007 8188 6071 8192
rect 6007 8132 6011 8188
rect 6011 8132 6067 8188
rect 6067 8132 6071 8188
rect 6007 8128 6071 8132
rect 6087 8188 6151 8192
rect 6087 8132 6091 8188
rect 6091 8132 6147 8188
rect 6147 8132 6151 8188
rect 6087 8128 6151 8132
rect 9111 8188 9175 8192
rect 9111 8132 9115 8188
rect 9115 8132 9171 8188
rect 9171 8132 9175 8188
rect 9111 8128 9175 8132
rect 9191 8188 9255 8192
rect 9191 8132 9195 8188
rect 9195 8132 9251 8188
rect 9251 8132 9255 8188
rect 9191 8128 9255 8132
rect 9271 8188 9335 8192
rect 9271 8132 9275 8188
rect 9275 8132 9331 8188
rect 9331 8132 9335 8188
rect 9271 8128 9335 8132
rect 9351 8188 9415 8192
rect 9351 8132 9355 8188
rect 9355 8132 9411 8188
rect 9411 8132 9415 8188
rect 9351 8128 9415 8132
rect 4215 7644 4279 7648
rect 4215 7588 4219 7644
rect 4219 7588 4275 7644
rect 4275 7588 4279 7644
rect 4215 7584 4279 7588
rect 4295 7644 4359 7648
rect 4295 7588 4299 7644
rect 4299 7588 4355 7644
rect 4355 7588 4359 7644
rect 4295 7584 4359 7588
rect 4375 7644 4439 7648
rect 4375 7588 4379 7644
rect 4379 7588 4435 7644
rect 4435 7588 4439 7644
rect 4375 7584 4439 7588
rect 4455 7644 4519 7648
rect 4455 7588 4459 7644
rect 4459 7588 4515 7644
rect 4515 7588 4519 7644
rect 4455 7584 4519 7588
rect 7479 7644 7543 7648
rect 7479 7588 7483 7644
rect 7483 7588 7539 7644
rect 7539 7588 7543 7644
rect 7479 7584 7543 7588
rect 7559 7644 7623 7648
rect 7559 7588 7563 7644
rect 7563 7588 7619 7644
rect 7619 7588 7623 7644
rect 7559 7584 7623 7588
rect 7639 7644 7703 7648
rect 7639 7588 7643 7644
rect 7643 7588 7699 7644
rect 7699 7588 7703 7644
rect 7639 7584 7703 7588
rect 7719 7644 7783 7648
rect 7719 7588 7723 7644
rect 7723 7588 7779 7644
rect 7779 7588 7783 7644
rect 7719 7584 7783 7588
rect 2584 7100 2648 7104
rect 2584 7044 2588 7100
rect 2588 7044 2644 7100
rect 2644 7044 2648 7100
rect 2584 7040 2648 7044
rect 2664 7100 2728 7104
rect 2664 7044 2668 7100
rect 2668 7044 2724 7100
rect 2724 7044 2728 7100
rect 2664 7040 2728 7044
rect 2744 7100 2808 7104
rect 2744 7044 2748 7100
rect 2748 7044 2804 7100
rect 2804 7044 2808 7100
rect 2744 7040 2808 7044
rect 2824 7100 2888 7104
rect 2824 7044 2828 7100
rect 2828 7044 2884 7100
rect 2884 7044 2888 7100
rect 2824 7040 2888 7044
rect 5847 7100 5911 7104
rect 5847 7044 5851 7100
rect 5851 7044 5907 7100
rect 5907 7044 5911 7100
rect 5847 7040 5911 7044
rect 5927 7100 5991 7104
rect 5927 7044 5931 7100
rect 5931 7044 5987 7100
rect 5987 7044 5991 7100
rect 5927 7040 5991 7044
rect 6007 7100 6071 7104
rect 6007 7044 6011 7100
rect 6011 7044 6067 7100
rect 6067 7044 6071 7100
rect 6007 7040 6071 7044
rect 6087 7100 6151 7104
rect 6087 7044 6091 7100
rect 6091 7044 6147 7100
rect 6147 7044 6151 7100
rect 6087 7040 6151 7044
rect 9111 7100 9175 7104
rect 9111 7044 9115 7100
rect 9115 7044 9171 7100
rect 9171 7044 9175 7100
rect 9111 7040 9175 7044
rect 9191 7100 9255 7104
rect 9191 7044 9195 7100
rect 9195 7044 9251 7100
rect 9251 7044 9255 7100
rect 9191 7040 9255 7044
rect 9271 7100 9335 7104
rect 9271 7044 9275 7100
rect 9275 7044 9331 7100
rect 9331 7044 9335 7100
rect 9271 7040 9335 7044
rect 9351 7100 9415 7104
rect 9351 7044 9355 7100
rect 9355 7044 9411 7100
rect 9411 7044 9415 7100
rect 9351 7040 9415 7044
rect 4215 6556 4279 6560
rect 4215 6500 4219 6556
rect 4219 6500 4275 6556
rect 4275 6500 4279 6556
rect 4215 6496 4279 6500
rect 4295 6556 4359 6560
rect 4295 6500 4299 6556
rect 4299 6500 4355 6556
rect 4355 6500 4359 6556
rect 4295 6496 4359 6500
rect 4375 6556 4439 6560
rect 4375 6500 4379 6556
rect 4379 6500 4435 6556
rect 4435 6500 4439 6556
rect 4375 6496 4439 6500
rect 4455 6556 4519 6560
rect 4455 6500 4459 6556
rect 4459 6500 4515 6556
rect 4515 6500 4519 6556
rect 4455 6496 4519 6500
rect 7479 6556 7543 6560
rect 7479 6500 7483 6556
rect 7483 6500 7539 6556
rect 7539 6500 7543 6556
rect 7479 6496 7543 6500
rect 7559 6556 7623 6560
rect 7559 6500 7563 6556
rect 7563 6500 7619 6556
rect 7619 6500 7623 6556
rect 7559 6496 7623 6500
rect 7639 6556 7703 6560
rect 7639 6500 7643 6556
rect 7643 6500 7699 6556
rect 7699 6500 7703 6556
rect 7639 6496 7703 6500
rect 7719 6556 7783 6560
rect 7719 6500 7723 6556
rect 7723 6500 7779 6556
rect 7779 6500 7783 6556
rect 7719 6496 7783 6500
rect 2584 6012 2648 6016
rect 2584 5956 2588 6012
rect 2588 5956 2644 6012
rect 2644 5956 2648 6012
rect 2584 5952 2648 5956
rect 2664 6012 2728 6016
rect 2664 5956 2668 6012
rect 2668 5956 2724 6012
rect 2724 5956 2728 6012
rect 2664 5952 2728 5956
rect 2744 6012 2808 6016
rect 2744 5956 2748 6012
rect 2748 5956 2804 6012
rect 2804 5956 2808 6012
rect 2744 5952 2808 5956
rect 2824 6012 2888 6016
rect 2824 5956 2828 6012
rect 2828 5956 2884 6012
rect 2884 5956 2888 6012
rect 2824 5952 2888 5956
rect 5847 6012 5911 6016
rect 5847 5956 5851 6012
rect 5851 5956 5907 6012
rect 5907 5956 5911 6012
rect 5847 5952 5911 5956
rect 5927 6012 5991 6016
rect 5927 5956 5931 6012
rect 5931 5956 5987 6012
rect 5987 5956 5991 6012
rect 5927 5952 5991 5956
rect 6007 6012 6071 6016
rect 6007 5956 6011 6012
rect 6011 5956 6067 6012
rect 6067 5956 6071 6012
rect 6007 5952 6071 5956
rect 6087 6012 6151 6016
rect 6087 5956 6091 6012
rect 6091 5956 6147 6012
rect 6147 5956 6151 6012
rect 6087 5952 6151 5956
rect 9111 6012 9175 6016
rect 9111 5956 9115 6012
rect 9115 5956 9171 6012
rect 9171 5956 9175 6012
rect 9111 5952 9175 5956
rect 9191 6012 9255 6016
rect 9191 5956 9195 6012
rect 9195 5956 9251 6012
rect 9251 5956 9255 6012
rect 9191 5952 9255 5956
rect 9271 6012 9335 6016
rect 9271 5956 9275 6012
rect 9275 5956 9331 6012
rect 9331 5956 9335 6012
rect 9271 5952 9335 5956
rect 9351 6012 9415 6016
rect 9351 5956 9355 6012
rect 9355 5956 9411 6012
rect 9411 5956 9415 6012
rect 9351 5952 9415 5956
rect 4215 5468 4279 5472
rect 4215 5412 4219 5468
rect 4219 5412 4275 5468
rect 4275 5412 4279 5468
rect 4215 5408 4279 5412
rect 4295 5468 4359 5472
rect 4295 5412 4299 5468
rect 4299 5412 4355 5468
rect 4355 5412 4359 5468
rect 4295 5408 4359 5412
rect 4375 5468 4439 5472
rect 4375 5412 4379 5468
rect 4379 5412 4435 5468
rect 4435 5412 4439 5468
rect 4375 5408 4439 5412
rect 4455 5468 4519 5472
rect 4455 5412 4459 5468
rect 4459 5412 4515 5468
rect 4515 5412 4519 5468
rect 4455 5408 4519 5412
rect 7479 5468 7543 5472
rect 7479 5412 7483 5468
rect 7483 5412 7539 5468
rect 7539 5412 7543 5468
rect 7479 5408 7543 5412
rect 7559 5468 7623 5472
rect 7559 5412 7563 5468
rect 7563 5412 7619 5468
rect 7619 5412 7623 5468
rect 7559 5408 7623 5412
rect 7639 5468 7703 5472
rect 7639 5412 7643 5468
rect 7643 5412 7699 5468
rect 7699 5412 7703 5468
rect 7639 5408 7703 5412
rect 7719 5468 7783 5472
rect 7719 5412 7723 5468
rect 7723 5412 7779 5468
rect 7779 5412 7783 5468
rect 7719 5408 7783 5412
rect 2584 4924 2648 4928
rect 2584 4868 2588 4924
rect 2588 4868 2644 4924
rect 2644 4868 2648 4924
rect 2584 4864 2648 4868
rect 2664 4924 2728 4928
rect 2664 4868 2668 4924
rect 2668 4868 2724 4924
rect 2724 4868 2728 4924
rect 2664 4864 2728 4868
rect 2744 4924 2808 4928
rect 2744 4868 2748 4924
rect 2748 4868 2804 4924
rect 2804 4868 2808 4924
rect 2744 4864 2808 4868
rect 2824 4924 2888 4928
rect 2824 4868 2828 4924
rect 2828 4868 2884 4924
rect 2884 4868 2888 4924
rect 2824 4864 2888 4868
rect 5847 4924 5911 4928
rect 5847 4868 5851 4924
rect 5851 4868 5907 4924
rect 5907 4868 5911 4924
rect 5847 4864 5911 4868
rect 5927 4924 5991 4928
rect 5927 4868 5931 4924
rect 5931 4868 5987 4924
rect 5987 4868 5991 4924
rect 5927 4864 5991 4868
rect 6007 4924 6071 4928
rect 6007 4868 6011 4924
rect 6011 4868 6067 4924
rect 6067 4868 6071 4924
rect 6007 4864 6071 4868
rect 6087 4924 6151 4928
rect 6087 4868 6091 4924
rect 6091 4868 6147 4924
rect 6147 4868 6151 4924
rect 6087 4864 6151 4868
rect 9111 4924 9175 4928
rect 9111 4868 9115 4924
rect 9115 4868 9171 4924
rect 9171 4868 9175 4924
rect 9111 4864 9175 4868
rect 9191 4924 9255 4928
rect 9191 4868 9195 4924
rect 9195 4868 9251 4924
rect 9251 4868 9255 4924
rect 9191 4864 9255 4868
rect 9271 4924 9335 4928
rect 9271 4868 9275 4924
rect 9275 4868 9331 4924
rect 9331 4868 9335 4924
rect 9271 4864 9335 4868
rect 9351 4924 9415 4928
rect 9351 4868 9355 4924
rect 9355 4868 9411 4924
rect 9411 4868 9415 4924
rect 9351 4864 9415 4868
rect 4215 4380 4279 4384
rect 4215 4324 4219 4380
rect 4219 4324 4275 4380
rect 4275 4324 4279 4380
rect 4215 4320 4279 4324
rect 4295 4380 4359 4384
rect 4295 4324 4299 4380
rect 4299 4324 4355 4380
rect 4355 4324 4359 4380
rect 4295 4320 4359 4324
rect 4375 4380 4439 4384
rect 4375 4324 4379 4380
rect 4379 4324 4435 4380
rect 4435 4324 4439 4380
rect 4375 4320 4439 4324
rect 4455 4380 4519 4384
rect 4455 4324 4459 4380
rect 4459 4324 4515 4380
rect 4515 4324 4519 4380
rect 4455 4320 4519 4324
rect 7479 4380 7543 4384
rect 7479 4324 7483 4380
rect 7483 4324 7539 4380
rect 7539 4324 7543 4380
rect 7479 4320 7543 4324
rect 7559 4380 7623 4384
rect 7559 4324 7563 4380
rect 7563 4324 7619 4380
rect 7619 4324 7623 4380
rect 7559 4320 7623 4324
rect 7639 4380 7703 4384
rect 7639 4324 7643 4380
rect 7643 4324 7699 4380
rect 7699 4324 7703 4380
rect 7639 4320 7703 4324
rect 7719 4380 7783 4384
rect 7719 4324 7723 4380
rect 7723 4324 7779 4380
rect 7779 4324 7783 4380
rect 7719 4320 7783 4324
rect 2584 3836 2648 3840
rect 2584 3780 2588 3836
rect 2588 3780 2644 3836
rect 2644 3780 2648 3836
rect 2584 3776 2648 3780
rect 2664 3836 2728 3840
rect 2664 3780 2668 3836
rect 2668 3780 2724 3836
rect 2724 3780 2728 3836
rect 2664 3776 2728 3780
rect 2744 3836 2808 3840
rect 2744 3780 2748 3836
rect 2748 3780 2804 3836
rect 2804 3780 2808 3836
rect 2744 3776 2808 3780
rect 2824 3836 2888 3840
rect 2824 3780 2828 3836
rect 2828 3780 2884 3836
rect 2884 3780 2888 3836
rect 2824 3776 2888 3780
rect 5847 3836 5911 3840
rect 5847 3780 5851 3836
rect 5851 3780 5907 3836
rect 5907 3780 5911 3836
rect 5847 3776 5911 3780
rect 5927 3836 5991 3840
rect 5927 3780 5931 3836
rect 5931 3780 5987 3836
rect 5987 3780 5991 3836
rect 5927 3776 5991 3780
rect 6007 3836 6071 3840
rect 6007 3780 6011 3836
rect 6011 3780 6067 3836
rect 6067 3780 6071 3836
rect 6007 3776 6071 3780
rect 6087 3836 6151 3840
rect 6087 3780 6091 3836
rect 6091 3780 6147 3836
rect 6147 3780 6151 3836
rect 6087 3776 6151 3780
rect 9111 3836 9175 3840
rect 9111 3780 9115 3836
rect 9115 3780 9171 3836
rect 9171 3780 9175 3836
rect 9111 3776 9175 3780
rect 9191 3836 9255 3840
rect 9191 3780 9195 3836
rect 9195 3780 9251 3836
rect 9251 3780 9255 3836
rect 9191 3776 9255 3780
rect 9271 3836 9335 3840
rect 9271 3780 9275 3836
rect 9275 3780 9331 3836
rect 9331 3780 9335 3836
rect 9271 3776 9335 3780
rect 9351 3836 9415 3840
rect 9351 3780 9355 3836
rect 9355 3780 9411 3836
rect 9411 3780 9415 3836
rect 9351 3776 9415 3780
rect 4215 3292 4279 3296
rect 4215 3236 4219 3292
rect 4219 3236 4275 3292
rect 4275 3236 4279 3292
rect 4215 3232 4279 3236
rect 4295 3292 4359 3296
rect 4295 3236 4299 3292
rect 4299 3236 4355 3292
rect 4355 3236 4359 3292
rect 4295 3232 4359 3236
rect 4375 3292 4439 3296
rect 4375 3236 4379 3292
rect 4379 3236 4435 3292
rect 4435 3236 4439 3292
rect 4375 3232 4439 3236
rect 4455 3292 4519 3296
rect 4455 3236 4459 3292
rect 4459 3236 4515 3292
rect 4515 3236 4519 3292
rect 4455 3232 4519 3236
rect 7479 3292 7543 3296
rect 7479 3236 7483 3292
rect 7483 3236 7539 3292
rect 7539 3236 7543 3292
rect 7479 3232 7543 3236
rect 7559 3292 7623 3296
rect 7559 3236 7563 3292
rect 7563 3236 7619 3292
rect 7619 3236 7623 3292
rect 7559 3232 7623 3236
rect 7639 3292 7703 3296
rect 7639 3236 7643 3292
rect 7643 3236 7699 3292
rect 7699 3236 7703 3292
rect 7639 3232 7703 3236
rect 7719 3292 7783 3296
rect 7719 3236 7723 3292
rect 7723 3236 7779 3292
rect 7779 3236 7783 3292
rect 7719 3232 7783 3236
rect 2584 2748 2648 2752
rect 2584 2692 2588 2748
rect 2588 2692 2644 2748
rect 2644 2692 2648 2748
rect 2584 2688 2648 2692
rect 2664 2748 2728 2752
rect 2664 2692 2668 2748
rect 2668 2692 2724 2748
rect 2724 2692 2728 2748
rect 2664 2688 2728 2692
rect 2744 2748 2808 2752
rect 2744 2692 2748 2748
rect 2748 2692 2804 2748
rect 2804 2692 2808 2748
rect 2744 2688 2808 2692
rect 2824 2748 2888 2752
rect 2824 2692 2828 2748
rect 2828 2692 2884 2748
rect 2884 2692 2888 2748
rect 2824 2688 2888 2692
rect 5847 2748 5911 2752
rect 5847 2692 5851 2748
rect 5851 2692 5907 2748
rect 5907 2692 5911 2748
rect 5847 2688 5911 2692
rect 5927 2748 5991 2752
rect 5927 2692 5931 2748
rect 5931 2692 5987 2748
rect 5987 2692 5991 2748
rect 5927 2688 5991 2692
rect 6007 2748 6071 2752
rect 6007 2692 6011 2748
rect 6011 2692 6067 2748
rect 6067 2692 6071 2748
rect 6007 2688 6071 2692
rect 6087 2748 6151 2752
rect 6087 2692 6091 2748
rect 6091 2692 6147 2748
rect 6147 2692 6151 2748
rect 6087 2688 6151 2692
rect 9111 2748 9175 2752
rect 9111 2692 9115 2748
rect 9115 2692 9171 2748
rect 9171 2692 9175 2748
rect 9111 2688 9175 2692
rect 9191 2748 9255 2752
rect 9191 2692 9195 2748
rect 9195 2692 9251 2748
rect 9251 2692 9255 2748
rect 9191 2688 9255 2692
rect 9271 2748 9335 2752
rect 9271 2692 9275 2748
rect 9275 2692 9331 2748
rect 9331 2692 9335 2748
rect 9271 2688 9335 2692
rect 9351 2748 9415 2752
rect 9351 2692 9355 2748
rect 9355 2692 9411 2748
rect 9411 2692 9415 2748
rect 9351 2688 9415 2692
rect 4215 2204 4279 2208
rect 4215 2148 4219 2204
rect 4219 2148 4275 2204
rect 4275 2148 4279 2204
rect 4215 2144 4279 2148
rect 4295 2204 4359 2208
rect 4295 2148 4299 2204
rect 4299 2148 4355 2204
rect 4355 2148 4359 2204
rect 4295 2144 4359 2148
rect 4375 2204 4439 2208
rect 4375 2148 4379 2204
rect 4379 2148 4435 2204
rect 4435 2148 4439 2204
rect 4375 2144 4439 2148
rect 4455 2204 4519 2208
rect 4455 2148 4459 2204
rect 4459 2148 4515 2204
rect 4515 2148 4519 2204
rect 4455 2144 4519 2148
rect 7479 2204 7543 2208
rect 7479 2148 7483 2204
rect 7483 2148 7539 2204
rect 7539 2148 7543 2204
rect 7479 2144 7543 2148
rect 7559 2204 7623 2208
rect 7559 2148 7563 2204
rect 7563 2148 7619 2204
rect 7619 2148 7623 2204
rect 7559 2144 7623 2148
rect 7639 2204 7703 2208
rect 7639 2148 7643 2204
rect 7643 2148 7699 2204
rect 7699 2148 7703 2204
rect 7639 2144 7703 2148
rect 7719 2204 7783 2208
rect 7719 2148 7723 2204
rect 7723 2148 7779 2204
rect 7779 2148 7783 2204
rect 7719 2144 7783 2148
<< metal4 >>
rect 2575 77824 2896 77840
rect 2575 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2575 76736 2896 77760
rect 2575 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2575 75648 2896 76672
rect 2575 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2575 74560 2896 75584
rect 2575 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2575 73472 2896 74496
rect 2575 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2575 72384 2896 73408
rect 2575 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2575 71296 2896 72320
rect 2575 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 1531 70548 1597 70549
rect 1531 70484 1532 70548
rect 1596 70484 1597 70548
rect 1531 70483 1597 70484
rect 1534 67829 1594 70483
rect 2575 70208 2896 71232
rect 2575 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2575 69120 2896 70144
rect 2575 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 1715 69052 1781 69053
rect 1715 68988 1716 69052
rect 1780 68988 1781 69052
rect 1715 68987 1781 68988
rect 1531 67828 1597 67829
rect 1531 67764 1532 67828
rect 1596 67764 1597 67828
rect 1531 67763 1597 67764
rect 1718 58309 1778 68987
rect 2083 68644 2149 68645
rect 2083 68580 2084 68644
rect 2148 68580 2149 68644
rect 2083 68579 2149 68580
rect 2086 62117 2146 68579
rect 2575 68032 2896 69056
rect 2575 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2575 66944 2896 67968
rect 2575 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2575 65856 2896 66880
rect 2575 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2267 64836 2333 64837
rect 2267 64772 2268 64836
rect 2332 64772 2333 64836
rect 2267 64771 2333 64772
rect 2083 62116 2149 62117
rect 2083 62052 2084 62116
rect 2148 62052 2149 62116
rect 2083 62051 2149 62052
rect 2270 61573 2330 64771
rect 2575 64768 2896 65792
rect 2575 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2575 63680 2896 64704
rect 2575 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2575 62592 2896 63616
rect 2575 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2267 61572 2333 61573
rect 2267 61508 2268 61572
rect 2332 61508 2333 61572
rect 2267 61507 2333 61508
rect 2575 61504 2896 62528
rect 2575 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2575 60416 2896 61440
rect 2575 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2575 59328 2896 60352
rect 2575 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 1715 58308 1781 58309
rect 1715 58244 1716 58308
rect 1780 58244 1781 58308
rect 1715 58243 1781 58244
rect 2575 58240 2896 59264
rect 2575 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2575 57152 2896 58176
rect 2575 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2575 56064 2896 57088
rect 4207 77280 4527 77840
rect 4207 77216 4215 77280
rect 4279 77216 4295 77280
rect 4359 77216 4375 77280
rect 4439 77216 4455 77280
rect 4519 77216 4527 77280
rect 4207 76192 4527 77216
rect 4207 76128 4215 76192
rect 4279 76128 4295 76192
rect 4359 76128 4375 76192
rect 4439 76128 4455 76192
rect 4519 76128 4527 76192
rect 4207 75104 4527 76128
rect 4207 75040 4215 75104
rect 4279 75040 4295 75104
rect 4359 75040 4375 75104
rect 4439 75040 4455 75104
rect 4519 75040 4527 75104
rect 4207 74016 4527 75040
rect 4207 73952 4215 74016
rect 4279 73952 4295 74016
rect 4359 73952 4375 74016
rect 4439 73952 4455 74016
rect 4519 73952 4527 74016
rect 4207 72928 4527 73952
rect 4207 72864 4215 72928
rect 4279 72864 4295 72928
rect 4359 72864 4375 72928
rect 4439 72864 4455 72928
rect 4519 72864 4527 72928
rect 4207 71840 4527 72864
rect 4207 71776 4215 71840
rect 4279 71776 4295 71840
rect 4359 71776 4375 71840
rect 4439 71776 4455 71840
rect 4519 71776 4527 71840
rect 4207 70752 4527 71776
rect 4207 70688 4215 70752
rect 4279 70688 4295 70752
rect 4359 70688 4375 70752
rect 4439 70688 4455 70752
rect 4519 70688 4527 70752
rect 4207 69664 4527 70688
rect 4207 69600 4215 69664
rect 4279 69600 4295 69664
rect 4359 69600 4375 69664
rect 4439 69600 4455 69664
rect 4519 69600 4527 69664
rect 4207 68576 4527 69600
rect 4207 68512 4215 68576
rect 4279 68512 4295 68576
rect 4359 68512 4375 68576
rect 4439 68512 4455 68576
rect 4519 68512 4527 68576
rect 4207 67488 4527 68512
rect 4207 67424 4215 67488
rect 4279 67424 4295 67488
rect 4359 67424 4375 67488
rect 4439 67424 4455 67488
rect 4519 67424 4527 67488
rect 4207 66400 4527 67424
rect 4207 66336 4215 66400
rect 4279 66336 4295 66400
rect 4359 66336 4375 66400
rect 4439 66336 4455 66400
rect 4519 66336 4527 66400
rect 4207 65312 4527 66336
rect 4207 65248 4215 65312
rect 4279 65248 4295 65312
rect 4359 65248 4375 65312
rect 4439 65248 4455 65312
rect 4519 65248 4527 65312
rect 4207 64224 4527 65248
rect 4207 64160 4215 64224
rect 4279 64160 4295 64224
rect 4359 64160 4375 64224
rect 4439 64160 4455 64224
rect 4519 64160 4527 64224
rect 4207 63136 4527 64160
rect 4207 63072 4215 63136
rect 4279 63072 4295 63136
rect 4359 63072 4375 63136
rect 4439 63072 4455 63136
rect 4519 63072 4527 63136
rect 4207 62048 4527 63072
rect 4207 61984 4215 62048
rect 4279 61984 4295 62048
rect 4359 61984 4375 62048
rect 4439 61984 4455 62048
rect 4519 61984 4527 62048
rect 4207 60960 4527 61984
rect 4207 60896 4215 60960
rect 4279 60896 4295 60960
rect 4359 60896 4375 60960
rect 4439 60896 4455 60960
rect 4519 60896 4527 60960
rect 4207 59872 4527 60896
rect 4207 59808 4215 59872
rect 4279 59808 4295 59872
rect 4359 59808 4375 59872
rect 4439 59808 4455 59872
rect 4519 59808 4527 59872
rect 4207 58784 4527 59808
rect 4207 58720 4215 58784
rect 4279 58720 4295 58784
rect 4359 58720 4375 58784
rect 4439 58720 4455 58784
rect 4519 58720 4527 58784
rect 4207 57696 4527 58720
rect 4207 57632 4215 57696
rect 4279 57632 4295 57696
rect 4359 57632 4375 57696
rect 4439 57632 4455 57696
rect 4519 57632 4527 57696
rect 3003 56676 3069 56677
rect 3003 56612 3004 56676
rect 3068 56612 3069 56676
rect 3003 56611 3069 56612
rect 2575 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 1163 55316 1229 55317
rect 1163 55252 1164 55316
rect 1228 55252 1229 55316
rect 1163 55251 1229 55252
rect 1166 23629 1226 55251
rect 2575 54976 2896 56000
rect 2575 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2575 53888 2896 54912
rect 2575 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2267 53412 2333 53413
rect 2267 53348 2268 53412
rect 2332 53348 2333 53412
rect 2267 53347 2333 53348
rect 2270 51237 2330 53347
rect 2575 52800 2896 53824
rect 2575 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2575 51712 2896 52736
rect 2575 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2267 51236 2333 51237
rect 2267 51172 2268 51236
rect 2332 51172 2333 51236
rect 2267 51171 2333 51172
rect 2575 50624 2896 51648
rect 2575 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2575 49536 2896 50560
rect 2575 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2575 48448 2896 49472
rect 2575 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2575 47360 2896 48384
rect 2575 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2575 46272 2896 47296
rect 3006 46885 3066 56611
rect 4207 56608 4527 57632
rect 4207 56544 4215 56608
rect 4279 56544 4295 56608
rect 4359 56544 4375 56608
rect 4439 56544 4455 56608
rect 4519 56544 4527 56608
rect 3187 55860 3253 55861
rect 3187 55796 3188 55860
rect 3252 55796 3253 55860
rect 3187 55795 3253 55796
rect 3190 50693 3250 55795
rect 4207 55520 4527 56544
rect 5839 77824 6159 77840
rect 5839 77760 5847 77824
rect 5911 77760 5927 77824
rect 5991 77760 6007 77824
rect 6071 77760 6087 77824
rect 6151 77760 6159 77824
rect 5839 76736 6159 77760
rect 5839 76672 5847 76736
rect 5911 76672 5927 76736
rect 5991 76672 6007 76736
rect 6071 76672 6087 76736
rect 6151 76672 6159 76736
rect 5839 75648 6159 76672
rect 5839 75584 5847 75648
rect 5911 75584 5927 75648
rect 5991 75584 6007 75648
rect 6071 75584 6087 75648
rect 6151 75584 6159 75648
rect 5839 74560 6159 75584
rect 5839 74496 5847 74560
rect 5911 74496 5927 74560
rect 5991 74496 6007 74560
rect 6071 74496 6087 74560
rect 6151 74496 6159 74560
rect 5839 73472 6159 74496
rect 5839 73408 5847 73472
rect 5911 73408 5927 73472
rect 5991 73408 6007 73472
rect 6071 73408 6087 73472
rect 6151 73408 6159 73472
rect 5839 72384 6159 73408
rect 5839 72320 5847 72384
rect 5911 72320 5927 72384
rect 5991 72320 6007 72384
rect 6071 72320 6087 72384
rect 6151 72320 6159 72384
rect 5839 71296 6159 72320
rect 5839 71232 5847 71296
rect 5911 71232 5927 71296
rect 5991 71232 6007 71296
rect 6071 71232 6087 71296
rect 6151 71232 6159 71296
rect 5839 70208 6159 71232
rect 5839 70144 5847 70208
rect 5911 70144 5927 70208
rect 5991 70144 6007 70208
rect 6071 70144 6087 70208
rect 6151 70144 6159 70208
rect 5839 69120 6159 70144
rect 5839 69056 5847 69120
rect 5911 69056 5927 69120
rect 5991 69056 6007 69120
rect 6071 69056 6087 69120
rect 6151 69056 6159 69120
rect 5839 68032 6159 69056
rect 5839 67968 5847 68032
rect 5911 67968 5927 68032
rect 5991 67968 6007 68032
rect 6071 67968 6087 68032
rect 6151 67968 6159 68032
rect 5839 66944 6159 67968
rect 5839 66880 5847 66944
rect 5911 66880 5927 66944
rect 5991 66880 6007 66944
rect 6071 66880 6087 66944
rect 6151 66880 6159 66944
rect 5839 65856 6159 66880
rect 5839 65792 5847 65856
rect 5911 65792 5927 65856
rect 5991 65792 6007 65856
rect 6071 65792 6087 65856
rect 6151 65792 6159 65856
rect 5839 64768 6159 65792
rect 5839 64704 5847 64768
rect 5911 64704 5927 64768
rect 5991 64704 6007 64768
rect 6071 64704 6087 64768
rect 6151 64704 6159 64768
rect 5839 63680 6159 64704
rect 5839 63616 5847 63680
rect 5911 63616 5927 63680
rect 5991 63616 6007 63680
rect 6071 63616 6087 63680
rect 6151 63616 6159 63680
rect 5839 62592 6159 63616
rect 5839 62528 5847 62592
rect 5911 62528 5927 62592
rect 5991 62528 6007 62592
rect 6071 62528 6087 62592
rect 6151 62528 6159 62592
rect 5839 61504 6159 62528
rect 5839 61440 5847 61504
rect 5911 61440 5927 61504
rect 5991 61440 6007 61504
rect 6071 61440 6087 61504
rect 6151 61440 6159 61504
rect 5839 60416 6159 61440
rect 5839 60352 5847 60416
rect 5911 60352 5927 60416
rect 5991 60352 6007 60416
rect 6071 60352 6087 60416
rect 6151 60352 6159 60416
rect 5839 59328 6159 60352
rect 5839 59264 5847 59328
rect 5911 59264 5927 59328
rect 5991 59264 6007 59328
rect 6071 59264 6087 59328
rect 6151 59264 6159 59328
rect 5839 58240 6159 59264
rect 5839 58176 5847 58240
rect 5911 58176 5927 58240
rect 5991 58176 6007 58240
rect 6071 58176 6087 58240
rect 6151 58176 6159 58240
rect 5839 57152 6159 58176
rect 5839 57088 5847 57152
rect 5911 57088 5927 57152
rect 5991 57088 6007 57152
rect 6071 57088 6087 57152
rect 6151 57088 6159 57152
rect 4659 56268 4725 56269
rect 4659 56204 4660 56268
rect 4724 56204 4725 56268
rect 4659 56203 4725 56204
rect 4207 55456 4215 55520
rect 4279 55456 4295 55520
rect 4359 55456 4375 55520
rect 4439 55456 4455 55520
rect 4519 55456 4527 55520
rect 3371 54772 3437 54773
rect 3371 54708 3372 54772
rect 3436 54708 3437 54772
rect 3371 54707 3437 54708
rect 3187 50692 3253 50693
rect 3187 50628 3188 50692
rect 3252 50628 3253 50692
rect 3187 50627 3253 50628
rect 3374 49333 3434 54707
rect 4207 54432 4527 55456
rect 4207 54368 4215 54432
rect 4279 54368 4295 54432
rect 4359 54368 4375 54432
rect 4439 54368 4455 54432
rect 4519 54368 4527 54432
rect 4207 53344 4527 54368
rect 4207 53280 4215 53344
rect 4279 53280 4295 53344
rect 4359 53280 4375 53344
rect 4439 53280 4455 53344
rect 4519 53280 4527 53344
rect 4207 52256 4527 53280
rect 4207 52192 4215 52256
rect 4279 52192 4295 52256
rect 4359 52192 4375 52256
rect 4439 52192 4455 52256
rect 4519 52192 4527 52256
rect 4207 51168 4527 52192
rect 4207 51104 4215 51168
rect 4279 51104 4295 51168
rect 4359 51104 4375 51168
rect 4439 51104 4455 51168
rect 4519 51104 4527 51168
rect 4207 50080 4527 51104
rect 4207 50016 4215 50080
rect 4279 50016 4295 50080
rect 4359 50016 4375 50080
rect 4439 50016 4455 50080
rect 4519 50016 4527 50080
rect 3371 49332 3437 49333
rect 3371 49268 3372 49332
rect 3436 49268 3437 49332
rect 3371 49267 3437 49268
rect 4207 48992 4527 50016
rect 4207 48928 4215 48992
rect 4279 48928 4295 48992
rect 4359 48928 4375 48992
rect 4439 48928 4455 48992
rect 4519 48928 4527 48992
rect 3739 48244 3805 48245
rect 3739 48180 3740 48244
rect 3804 48180 3805 48244
rect 3739 48179 3805 48180
rect 3003 46884 3069 46885
rect 3003 46820 3004 46884
rect 3068 46820 3069 46884
rect 3003 46819 3069 46820
rect 2575 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2267 46068 2333 46069
rect 2267 46004 2268 46068
rect 2332 46004 2333 46068
rect 2267 46003 2333 46004
rect 2083 40356 2149 40357
rect 2083 40292 2084 40356
rect 2148 40292 2149 40356
rect 2083 40291 2149 40292
rect 2086 36821 2146 40291
rect 2270 40085 2330 46003
rect 2575 45184 2896 46208
rect 2575 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2575 44096 2896 45120
rect 2575 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2575 43008 2896 44032
rect 3742 43213 3802 48179
rect 4207 47904 4527 48928
rect 4662 48789 4722 56203
rect 5839 56064 6159 57088
rect 5839 56000 5847 56064
rect 5911 56000 5927 56064
rect 5991 56000 6007 56064
rect 6071 56000 6087 56064
rect 6151 56000 6159 56064
rect 5839 54976 6159 56000
rect 5839 54912 5847 54976
rect 5911 54912 5927 54976
rect 5991 54912 6007 54976
rect 6071 54912 6087 54976
rect 6151 54912 6159 54976
rect 5839 53888 6159 54912
rect 5839 53824 5847 53888
rect 5911 53824 5927 53888
rect 5991 53824 6007 53888
rect 6071 53824 6087 53888
rect 6151 53824 6159 53888
rect 5395 53684 5461 53685
rect 5395 53620 5396 53684
rect 5460 53620 5461 53684
rect 5395 53619 5461 53620
rect 4843 53140 4909 53141
rect 4843 53076 4844 53140
rect 4908 53076 4909 53140
rect 4843 53075 4909 53076
rect 4846 51645 4906 53075
rect 4843 51644 4909 51645
rect 4843 51580 4844 51644
rect 4908 51580 4909 51644
rect 4843 51579 4909 51580
rect 5398 51101 5458 53619
rect 5839 52800 6159 53824
rect 5839 52736 5847 52800
rect 5911 52736 5927 52800
rect 5991 52736 6007 52800
rect 6071 52736 6087 52800
rect 6151 52736 6159 52800
rect 5839 51712 6159 52736
rect 5839 51648 5847 51712
rect 5911 51648 5927 51712
rect 5991 51648 6007 51712
rect 6071 51648 6087 51712
rect 6151 51648 6159 51712
rect 5395 51100 5461 51101
rect 5395 51036 5396 51100
rect 5460 51036 5461 51100
rect 5395 51035 5461 51036
rect 5839 50624 6159 51648
rect 5839 50560 5847 50624
rect 5911 50560 5927 50624
rect 5991 50560 6007 50624
rect 6071 50560 6087 50624
rect 6151 50560 6159 50624
rect 5839 49536 6159 50560
rect 5839 49472 5847 49536
rect 5911 49472 5927 49536
rect 5991 49472 6007 49536
rect 6071 49472 6087 49536
rect 6151 49472 6159 49536
rect 4659 48788 4725 48789
rect 4659 48724 4660 48788
rect 4724 48724 4725 48788
rect 4659 48723 4725 48724
rect 5839 48448 6159 49472
rect 7471 77280 7791 77840
rect 7471 77216 7479 77280
rect 7543 77216 7559 77280
rect 7623 77216 7639 77280
rect 7703 77216 7719 77280
rect 7783 77216 7791 77280
rect 7471 76192 7791 77216
rect 7471 76128 7479 76192
rect 7543 76128 7559 76192
rect 7623 76128 7639 76192
rect 7703 76128 7719 76192
rect 7783 76128 7791 76192
rect 7471 75104 7791 76128
rect 7471 75040 7479 75104
rect 7543 75040 7559 75104
rect 7623 75040 7639 75104
rect 7703 75040 7719 75104
rect 7783 75040 7791 75104
rect 7471 74016 7791 75040
rect 7471 73952 7479 74016
rect 7543 73952 7559 74016
rect 7623 73952 7639 74016
rect 7703 73952 7719 74016
rect 7783 73952 7791 74016
rect 7471 72928 7791 73952
rect 7471 72864 7479 72928
rect 7543 72864 7559 72928
rect 7623 72864 7639 72928
rect 7703 72864 7719 72928
rect 7783 72864 7791 72928
rect 7471 71840 7791 72864
rect 7471 71776 7479 71840
rect 7543 71776 7559 71840
rect 7623 71776 7639 71840
rect 7703 71776 7719 71840
rect 7783 71776 7791 71840
rect 7471 70752 7791 71776
rect 7471 70688 7479 70752
rect 7543 70688 7559 70752
rect 7623 70688 7639 70752
rect 7703 70688 7719 70752
rect 7783 70688 7791 70752
rect 7471 69664 7791 70688
rect 7471 69600 7479 69664
rect 7543 69600 7559 69664
rect 7623 69600 7639 69664
rect 7703 69600 7719 69664
rect 7783 69600 7791 69664
rect 7471 68576 7791 69600
rect 7471 68512 7479 68576
rect 7543 68512 7559 68576
rect 7623 68512 7639 68576
rect 7703 68512 7719 68576
rect 7783 68512 7791 68576
rect 7471 67488 7791 68512
rect 7471 67424 7479 67488
rect 7543 67424 7559 67488
rect 7623 67424 7639 67488
rect 7703 67424 7719 67488
rect 7783 67424 7791 67488
rect 7471 66400 7791 67424
rect 7471 66336 7479 66400
rect 7543 66336 7559 66400
rect 7623 66336 7639 66400
rect 7703 66336 7719 66400
rect 7783 66336 7791 66400
rect 7471 65312 7791 66336
rect 7471 65248 7479 65312
rect 7543 65248 7559 65312
rect 7623 65248 7639 65312
rect 7703 65248 7719 65312
rect 7783 65248 7791 65312
rect 7471 64224 7791 65248
rect 7471 64160 7479 64224
rect 7543 64160 7559 64224
rect 7623 64160 7639 64224
rect 7703 64160 7719 64224
rect 7783 64160 7791 64224
rect 7471 63136 7791 64160
rect 7471 63072 7479 63136
rect 7543 63072 7559 63136
rect 7623 63072 7639 63136
rect 7703 63072 7719 63136
rect 7783 63072 7791 63136
rect 7471 62048 7791 63072
rect 7471 61984 7479 62048
rect 7543 61984 7559 62048
rect 7623 61984 7639 62048
rect 7703 61984 7719 62048
rect 7783 61984 7791 62048
rect 7471 60960 7791 61984
rect 7471 60896 7479 60960
rect 7543 60896 7559 60960
rect 7623 60896 7639 60960
rect 7703 60896 7719 60960
rect 7783 60896 7791 60960
rect 7471 59872 7791 60896
rect 7471 59808 7479 59872
rect 7543 59808 7559 59872
rect 7623 59808 7639 59872
rect 7703 59808 7719 59872
rect 7783 59808 7791 59872
rect 7471 58784 7791 59808
rect 7471 58720 7479 58784
rect 7543 58720 7559 58784
rect 7623 58720 7639 58784
rect 7703 58720 7719 58784
rect 7783 58720 7791 58784
rect 7471 57696 7791 58720
rect 7471 57632 7479 57696
rect 7543 57632 7559 57696
rect 7623 57632 7639 57696
rect 7703 57632 7719 57696
rect 7783 57632 7791 57696
rect 7471 56608 7791 57632
rect 7471 56544 7479 56608
rect 7543 56544 7559 56608
rect 7623 56544 7639 56608
rect 7703 56544 7719 56608
rect 7783 56544 7791 56608
rect 7471 55520 7791 56544
rect 7471 55456 7479 55520
rect 7543 55456 7559 55520
rect 7623 55456 7639 55520
rect 7703 55456 7719 55520
rect 7783 55456 7791 55520
rect 7471 54432 7791 55456
rect 7471 54368 7479 54432
rect 7543 54368 7559 54432
rect 7623 54368 7639 54432
rect 7703 54368 7719 54432
rect 7783 54368 7791 54432
rect 7471 53344 7791 54368
rect 7471 53280 7479 53344
rect 7543 53280 7559 53344
rect 7623 53280 7639 53344
rect 7703 53280 7719 53344
rect 7783 53280 7791 53344
rect 7471 52256 7791 53280
rect 7471 52192 7479 52256
rect 7543 52192 7559 52256
rect 7623 52192 7639 52256
rect 7703 52192 7719 52256
rect 7783 52192 7791 52256
rect 7471 51168 7791 52192
rect 7471 51104 7479 51168
rect 7543 51104 7559 51168
rect 7623 51104 7639 51168
rect 7703 51104 7719 51168
rect 7783 51104 7791 51168
rect 7471 50080 7791 51104
rect 7471 50016 7479 50080
rect 7543 50016 7559 50080
rect 7623 50016 7639 50080
rect 7703 50016 7719 50080
rect 7783 50016 7791 50080
rect 7471 48992 7791 50016
rect 7471 48928 7479 48992
rect 7543 48928 7559 48992
rect 7623 48928 7639 48992
rect 7703 48928 7719 48992
rect 7783 48928 7791 48992
rect 6683 48788 6749 48789
rect 6683 48724 6684 48788
rect 6748 48724 6749 48788
rect 6683 48723 6749 48724
rect 5839 48384 5847 48448
rect 5911 48384 5927 48448
rect 5991 48384 6007 48448
rect 6071 48384 6087 48448
rect 6151 48384 6159 48448
rect 4659 48108 4725 48109
rect 4659 48044 4660 48108
rect 4724 48044 4725 48108
rect 4659 48043 4725 48044
rect 4207 47840 4215 47904
rect 4279 47840 4295 47904
rect 4359 47840 4375 47904
rect 4439 47840 4455 47904
rect 4519 47840 4527 47904
rect 4207 46816 4527 47840
rect 4207 46752 4215 46816
rect 4279 46752 4295 46816
rect 4359 46752 4375 46816
rect 4439 46752 4455 46816
rect 4519 46752 4527 46816
rect 4207 45728 4527 46752
rect 4207 45664 4215 45728
rect 4279 45664 4295 45728
rect 4359 45664 4375 45728
rect 4439 45664 4455 45728
rect 4519 45664 4527 45728
rect 4207 44640 4527 45664
rect 4207 44576 4215 44640
rect 4279 44576 4295 44640
rect 4359 44576 4375 44640
rect 4439 44576 4455 44640
rect 4519 44576 4527 44640
rect 4207 43552 4527 44576
rect 4207 43488 4215 43552
rect 4279 43488 4295 43552
rect 4359 43488 4375 43552
rect 4439 43488 4455 43552
rect 4519 43488 4527 43552
rect 3739 43212 3805 43213
rect 3739 43148 3740 43212
rect 3804 43148 3805 43212
rect 3739 43147 3805 43148
rect 2575 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2575 41920 2896 42944
rect 2575 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2575 40832 2896 41856
rect 2575 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2267 40084 2333 40085
rect 2267 40020 2268 40084
rect 2332 40020 2333 40084
rect 2267 40019 2333 40020
rect 2575 39744 2896 40768
rect 2575 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2575 38656 2896 39680
rect 2575 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2575 37568 2896 38592
rect 2575 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2083 36820 2149 36821
rect 2083 36756 2084 36820
rect 2148 36756 2149 36820
rect 2083 36755 2149 36756
rect 2575 36480 2896 37504
rect 2575 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2575 35392 2896 36416
rect 2575 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2575 34304 2896 35328
rect 2575 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2575 33216 2896 34240
rect 2575 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2575 32128 2896 33152
rect 2575 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2575 31040 2896 32064
rect 2575 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2575 29952 2896 30976
rect 2575 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2575 28864 2896 29888
rect 2575 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2575 27776 2896 28800
rect 2575 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2575 26688 2896 27712
rect 2575 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2575 25600 2896 26624
rect 2575 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2575 24512 2896 25536
rect 2575 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 1163 23628 1229 23629
rect 1163 23564 1164 23628
rect 1228 23564 1229 23628
rect 1163 23563 1229 23564
rect 2575 23424 2896 24448
rect 2575 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2575 22336 2896 23360
rect 2575 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2575 21248 2896 22272
rect 2575 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2575 20160 2896 21184
rect 2575 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2575 19072 2896 20096
rect 2575 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2575 17984 2896 19008
rect 2575 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2575 16896 2896 17920
rect 2575 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2575 15808 2896 16832
rect 2575 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2575 14720 2896 15744
rect 2575 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2575 13632 2896 14656
rect 2575 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2575 12544 2896 13568
rect 2575 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2575 11456 2896 12480
rect 2575 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2575 10368 2896 11392
rect 2575 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2575 9280 2896 10304
rect 2575 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2575 8192 2896 9216
rect 2575 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2575 7104 2896 8128
rect 2575 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2575 6016 2896 7040
rect 2575 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2575 4928 2896 5952
rect 2575 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2575 3840 2896 4864
rect 2575 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2575 2752 2896 3776
rect 2575 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2575 2128 2896 2688
rect 4207 42464 4527 43488
rect 4207 42400 4215 42464
rect 4279 42400 4295 42464
rect 4359 42400 4375 42464
rect 4439 42400 4455 42464
rect 4519 42400 4527 42464
rect 4207 41376 4527 42400
rect 4662 41445 4722 48043
rect 5839 47360 6159 48384
rect 5839 47296 5847 47360
rect 5911 47296 5927 47360
rect 5991 47296 6007 47360
rect 6071 47296 6087 47360
rect 6151 47296 6159 47360
rect 5839 46272 6159 47296
rect 6686 46341 6746 48723
rect 7471 47904 7791 48928
rect 7471 47840 7479 47904
rect 7543 47840 7559 47904
rect 7623 47840 7639 47904
rect 7703 47840 7719 47904
rect 7783 47840 7791 47904
rect 7471 46816 7791 47840
rect 7471 46752 7479 46816
rect 7543 46752 7559 46816
rect 7623 46752 7639 46816
rect 7703 46752 7719 46816
rect 7783 46752 7791 46816
rect 6683 46340 6749 46341
rect 6683 46276 6684 46340
rect 6748 46276 6749 46340
rect 6683 46275 6749 46276
rect 5839 46208 5847 46272
rect 5911 46208 5927 46272
rect 5991 46208 6007 46272
rect 6071 46208 6087 46272
rect 6151 46208 6159 46272
rect 5839 45184 6159 46208
rect 5839 45120 5847 45184
rect 5911 45120 5927 45184
rect 5991 45120 6007 45184
rect 6071 45120 6087 45184
rect 6151 45120 6159 45184
rect 5839 44096 6159 45120
rect 5839 44032 5847 44096
rect 5911 44032 5927 44096
rect 5991 44032 6007 44096
rect 6071 44032 6087 44096
rect 6151 44032 6159 44096
rect 5839 43008 6159 44032
rect 5839 42944 5847 43008
rect 5911 42944 5927 43008
rect 5991 42944 6007 43008
rect 6071 42944 6087 43008
rect 6151 42944 6159 43008
rect 5839 41920 6159 42944
rect 5839 41856 5847 41920
rect 5911 41856 5927 41920
rect 5991 41856 6007 41920
rect 6071 41856 6087 41920
rect 6151 41856 6159 41920
rect 4659 41444 4725 41445
rect 4659 41380 4660 41444
rect 4724 41380 4725 41444
rect 4659 41379 4725 41380
rect 4207 41312 4215 41376
rect 4279 41312 4295 41376
rect 4359 41312 4375 41376
rect 4439 41312 4455 41376
rect 4519 41312 4527 41376
rect 4207 40288 4527 41312
rect 4207 40224 4215 40288
rect 4279 40224 4295 40288
rect 4359 40224 4375 40288
rect 4439 40224 4455 40288
rect 4519 40224 4527 40288
rect 4207 39200 4527 40224
rect 4207 39136 4215 39200
rect 4279 39136 4295 39200
rect 4359 39136 4375 39200
rect 4439 39136 4455 39200
rect 4519 39136 4527 39200
rect 4207 38112 4527 39136
rect 4207 38048 4215 38112
rect 4279 38048 4295 38112
rect 4359 38048 4375 38112
rect 4439 38048 4455 38112
rect 4519 38048 4527 38112
rect 4207 37024 4527 38048
rect 4207 36960 4215 37024
rect 4279 36960 4295 37024
rect 4359 36960 4375 37024
rect 4439 36960 4455 37024
rect 4519 36960 4527 37024
rect 4207 35936 4527 36960
rect 4207 35872 4215 35936
rect 4279 35872 4295 35936
rect 4359 35872 4375 35936
rect 4439 35872 4455 35936
rect 4519 35872 4527 35936
rect 4207 34848 4527 35872
rect 4207 34784 4215 34848
rect 4279 34784 4295 34848
rect 4359 34784 4375 34848
rect 4439 34784 4455 34848
rect 4519 34784 4527 34848
rect 4207 33760 4527 34784
rect 4207 33696 4215 33760
rect 4279 33696 4295 33760
rect 4359 33696 4375 33760
rect 4439 33696 4455 33760
rect 4519 33696 4527 33760
rect 4207 32672 4527 33696
rect 4207 32608 4215 32672
rect 4279 32608 4295 32672
rect 4359 32608 4375 32672
rect 4439 32608 4455 32672
rect 4519 32608 4527 32672
rect 4207 31584 4527 32608
rect 4207 31520 4215 31584
rect 4279 31520 4295 31584
rect 4359 31520 4375 31584
rect 4439 31520 4455 31584
rect 4519 31520 4527 31584
rect 4207 30496 4527 31520
rect 4207 30432 4215 30496
rect 4279 30432 4295 30496
rect 4359 30432 4375 30496
rect 4439 30432 4455 30496
rect 4519 30432 4527 30496
rect 4207 29408 4527 30432
rect 4207 29344 4215 29408
rect 4279 29344 4295 29408
rect 4359 29344 4375 29408
rect 4439 29344 4455 29408
rect 4519 29344 4527 29408
rect 4207 28320 4527 29344
rect 4207 28256 4215 28320
rect 4279 28256 4295 28320
rect 4359 28256 4375 28320
rect 4439 28256 4455 28320
rect 4519 28256 4527 28320
rect 4207 27232 4527 28256
rect 4207 27168 4215 27232
rect 4279 27168 4295 27232
rect 4359 27168 4375 27232
rect 4439 27168 4455 27232
rect 4519 27168 4527 27232
rect 4207 26144 4527 27168
rect 4207 26080 4215 26144
rect 4279 26080 4295 26144
rect 4359 26080 4375 26144
rect 4439 26080 4455 26144
rect 4519 26080 4527 26144
rect 4207 25056 4527 26080
rect 4207 24992 4215 25056
rect 4279 24992 4295 25056
rect 4359 24992 4375 25056
rect 4439 24992 4455 25056
rect 4519 24992 4527 25056
rect 4207 23968 4527 24992
rect 4207 23904 4215 23968
rect 4279 23904 4295 23968
rect 4359 23904 4375 23968
rect 4439 23904 4455 23968
rect 4519 23904 4527 23968
rect 4207 22880 4527 23904
rect 4207 22816 4215 22880
rect 4279 22816 4295 22880
rect 4359 22816 4375 22880
rect 4439 22816 4455 22880
rect 4519 22816 4527 22880
rect 4207 21792 4527 22816
rect 4207 21728 4215 21792
rect 4279 21728 4295 21792
rect 4359 21728 4375 21792
rect 4439 21728 4455 21792
rect 4519 21728 4527 21792
rect 4207 20704 4527 21728
rect 4207 20640 4215 20704
rect 4279 20640 4295 20704
rect 4359 20640 4375 20704
rect 4439 20640 4455 20704
rect 4519 20640 4527 20704
rect 4207 19616 4527 20640
rect 4207 19552 4215 19616
rect 4279 19552 4295 19616
rect 4359 19552 4375 19616
rect 4439 19552 4455 19616
rect 4519 19552 4527 19616
rect 4207 18528 4527 19552
rect 4207 18464 4215 18528
rect 4279 18464 4295 18528
rect 4359 18464 4375 18528
rect 4439 18464 4455 18528
rect 4519 18464 4527 18528
rect 4207 17440 4527 18464
rect 4207 17376 4215 17440
rect 4279 17376 4295 17440
rect 4359 17376 4375 17440
rect 4439 17376 4455 17440
rect 4519 17376 4527 17440
rect 4207 16352 4527 17376
rect 4207 16288 4215 16352
rect 4279 16288 4295 16352
rect 4359 16288 4375 16352
rect 4439 16288 4455 16352
rect 4519 16288 4527 16352
rect 4207 15264 4527 16288
rect 4207 15200 4215 15264
rect 4279 15200 4295 15264
rect 4359 15200 4375 15264
rect 4439 15200 4455 15264
rect 4519 15200 4527 15264
rect 4207 14176 4527 15200
rect 4207 14112 4215 14176
rect 4279 14112 4295 14176
rect 4359 14112 4375 14176
rect 4439 14112 4455 14176
rect 4519 14112 4527 14176
rect 4207 13088 4527 14112
rect 4207 13024 4215 13088
rect 4279 13024 4295 13088
rect 4359 13024 4375 13088
rect 4439 13024 4455 13088
rect 4519 13024 4527 13088
rect 4207 12000 4527 13024
rect 4207 11936 4215 12000
rect 4279 11936 4295 12000
rect 4359 11936 4375 12000
rect 4439 11936 4455 12000
rect 4519 11936 4527 12000
rect 4207 10912 4527 11936
rect 4207 10848 4215 10912
rect 4279 10848 4295 10912
rect 4359 10848 4375 10912
rect 4439 10848 4455 10912
rect 4519 10848 4527 10912
rect 4207 9824 4527 10848
rect 4207 9760 4215 9824
rect 4279 9760 4295 9824
rect 4359 9760 4375 9824
rect 4439 9760 4455 9824
rect 4519 9760 4527 9824
rect 4207 8736 4527 9760
rect 4207 8672 4215 8736
rect 4279 8672 4295 8736
rect 4359 8672 4375 8736
rect 4439 8672 4455 8736
rect 4519 8672 4527 8736
rect 4207 7648 4527 8672
rect 4207 7584 4215 7648
rect 4279 7584 4295 7648
rect 4359 7584 4375 7648
rect 4439 7584 4455 7648
rect 4519 7584 4527 7648
rect 4207 6560 4527 7584
rect 4207 6496 4215 6560
rect 4279 6496 4295 6560
rect 4359 6496 4375 6560
rect 4439 6496 4455 6560
rect 4519 6496 4527 6560
rect 4207 5472 4527 6496
rect 4207 5408 4215 5472
rect 4279 5408 4295 5472
rect 4359 5408 4375 5472
rect 4439 5408 4455 5472
rect 4519 5408 4527 5472
rect 4207 4384 4527 5408
rect 4207 4320 4215 4384
rect 4279 4320 4295 4384
rect 4359 4320 4375 4384
rect 4439 4320 4455 4384
rect 4519 4320 4527 4384
rect 4207 3296 4527 4320
rect 4207 3232 4215 3296
rect 4279 3232 4295 3296
rect 4359 3232 4375 3296
rect 4439 3232 4455 3296
rect 4519 3232 4527 3296
rect 4207 2208 4527 3232
rect 4207 2144 4215 2208
rect 4279 2144 4295 2208
rect 4359 2144 4375 2208
rect 4439 2144 4455 2208
rect 4519 2144 4527 2208
rect 4207 2128 4527 2144
rect 5839 40832 6159 41856
rect 5839 40768 5847 40832
rect 5911 40768 5927 40832
rect 5991 40768 6007 40832
rect 6071 40768 6087 40832
rect 6151 40768 6159 40832
rect 5839 39744 6159 40768
rect 5839 39680 5847 39744
rect 5911 39680 5927 39744
rect 5991 39680 6007 39744
rect 6071 39680 6087 39744
rect 6151 39680 6159 39744
rect 5839 38656 6159 39680
rect 5839 38592 5847 38656
rect 5911 38592 5927 38656
rect 5991 38592 6007 38656
rect 6071 38592 6087 38656
rect 6151 38592 6159 38656
rect 5839 37568 6159 38592
rect 5839 37504 5847 37568
rect 5911 37504 5927 37568
rect 5991 37504 6007 37568
rect 6071 37504 6087 37568
rect 6151 37504 6159 37568
rect 5839 36480 6159 37504
rect 5839 36416 5847 36480
rect 5911 36416 5927 36480
rect 5991 36416 6007 36480
rect 6071 36416 6087 36480
rect 6151 36416 6159 36480
rect 5839 35392 6159 36416
rect 5839 35328 5847 35392
rect 5911 35328 5927 35392
rect 5991 35328 6007 35392
rect 6071 35328 6087 35392
rect 6151 35328 6159 35392
rect 5839 34304 6159 35328
rect 5839 34240 5847 34304
rect 5911 34240 5927 34304
rect 5991 34240 6007 34304
rect 6071 34240 6087 34304
rect 6151 34240 6159 34304
rect 5839 33216 6159 34240
rect 5839 33152 5847 33216
rect 5911 33152 5927 33216
rect 5991 33152 6007 33216
rect 6071 33152 6087 33216
rect 6151 33152 6159 33216
rect 5839 32128 6159 33152
rect 5839 32064 5847 32128
rect 5911 32064 5927 32128
rect 5991 32064 6007 32128
rect 6071 32064 6087 32128
rect 6151 32064 6159 32128
rect 5839 31040 6159 32064
rect 5839 30976 5847 31040
rect 5911 30976 5927 31040
rect 5991 30976 6007 31040
rect 6071 30976 6087 31040
rect 6151 30976 6159 31040
rect 5839 29952 6159 30976
rect 5839 29888 5847 29952
rect 5911 29888 5927 29952
rect 5991 29888 6007 29952
rect 6071 29888 6087 29952
rect 6151 29888 6159 29952
rect 5839 28864 6159 29888
rect 5839 28800 5847 28864
rect 5911 28800 5927 28864
rect 5991 28800 6007 28864
rect 6071 28800 6087 28864
rect 6151 28800 6159 28864
rect 5839 27776 6159 28800
rect 5839 27712 5847 27776
rect 5911 27712 5927 27776
rect 5991 27712 6007 27776
rect 6071 27712 6087 27776
rect 6151 27712 6159 27776
rect 5839 26688 6159 27712
rect 5839 26624 5847 26688
rect 5911 26624 5927 26688
rect 5991 26624 6007 26688
rect 6071 26624 6087 26688
rect 6151 26624 6159 26688
rect 5839 25600 6159 26624
rect 5839 25536 5847 25600
rect 5911 25536 5927 25600
rect 5991 25536 6007 25600
rect 6071 25536 6087 25600
rect 6151 25536 6159 25600
rect 5839 24512 6159 25536
rect 5839 24448 5847 24512
rect 5911 24448 5927 24512
rect 5991 24448 6007 24512
rect 6071 24448 6087 24512
rect 6151 24448 6159 24512
rect 5839 23424 6159 24448
rect 5839 23360 5847 23424
rect 5911 23360 5927 23424
rect 5991 23360 6007 23424
rect 6071 23360 6087 23424
rect 6151 23360 6159 23424
rect 5839 22336 6159 23360
rect 5839 22272 5847 22336
rect 5911 22272 5927 22336
rect 5991 22272 6007 22336
rect 6071 22272 6087 22336
rect 6151 22272 6159 22336
rect 5839 21248 6159 22272
rect 5839 21184 5847 21248
rect 5911 21184 5927 21248
rect 5991 21184 6007 21248
rect 6071 21184 6087 21248
rect 6151 21184 6159 21248
rect 5839 20160 6159 21184
rect 5839 20096 5847 20160
rect 5911 20096 5927 20160
rect 5991 20096 6007 20160
rect 6071 20096 6087 20160
rect 6151 20096 6159 20160
rect 5839 19072 6159 20096
rect 5839 19008 5847 19072
rect 5911 19008 5927 19072
rect 5991 19008 6007 19072
rect 6071 19008 6087 19072
rect 6151 19008 6159 19072
rect 5839 17984 6159 19008
rect 5839 17920 5847 17984
rect 5911 17920 5927 17984
rect 5991 17920 6007 17984
rect 6071 17920 6087 17984
rect 6151 17920 6159 17984
rect 5839 16896 6159 17920
rect 5839 16832 5847 16896
rect 5911 16832 5927 16896
rect 5991 16832 6007 16896
rect 6071 16832 6087 16896
rect 6151 16832 6159 16896
rect 5839 15808 6159 16832
rect 5839 15744 5847 15808
rect 5911 15744 5927 15808
rect 5991 15744 6007 15808
rect 6071 15744 6087 15808
rect 6151 15744 6159 15808
rect 5839 14720 6159 15744
rect 5839 14656 5847 14720
rect 5911 14656 5927 14720
rect 5991 14656 6007 14720
rect 6071 14656 6087 14720
rect 6151 14656 6159 14720
rect 5839 13632 6159 14656
rect 5839 13568 5847 13632
rect 5911 13568 5927 13632
rect 5991 13568 6007 13632
rect 6071 13568 6087 13632
rect 6151 13568 6159 13632
rect 5839 12544 6159 13568
rect 5839 12480 5847 12544
rect 5911 12480 5927 12544
rect 5991 12480 6007 12544
rect 6071 12480 6087 12544
rect 6151 12480 6159 12544
rect 5839 11456 6159 12480
rect 5839 11392 5847 11456
rect 5911 11392 5927 11456
rect 5991 11392 6007 11456
rect 6071 11392 6087 11456
rect 6151 11392 6159 11456
rect 5839 10368 6159 11392
rect 5839 10304 5847 10368
rect 5911 10304 5927 10368
rect 5991 10304 6007 10368
rect 6071 10304 6087 10368
rect 6151 10304 6159 10368
rect 5839 9280 6159 10304
rect 5839 9216 5847 9280
rect 5911 9216 5927 9280
rect 5991 9216 6007 9280
rect 6071 9216 6087 9280
rect 6151 9216 6159 9280
rect 5839 8192 6159 9216
rect 5839 8128 5847 8192
rect 5911 8128 5927 8192
rect 5991 8128 6007 8192
rect 6071 8128 6087 8192
rect 6151 8128 6159 8192
rect 5839 7104 6159 8128
rect 5839 7040 5847 7104
rect 5911 7040 5927 7104
rect 5991 7040 6007 7104
rect 6071 7040 6087 7104
rect 6151 7040 6159 7104
rect 5839 6016 6159 7040
rect 5839 5952 5847 6016
rect 5911 5952 5927 6016
rect 5991 5952 6007 6016
rect 6071 5952 6087 6016
rect 6151 5952 6159 6016
rect 5839 4928 6159 5952
rect 5839 4864 5847 4928
rect 5911 4864 5927 4928
rect 5991 4864 6007 4928
rect 6071 4864 6087 4928
rect 6151 4864 6159 4928
rect 5839 3840 6159 4864
rect 5839 3776 5847 3840
rect 5911 3776 5927 3840
rect 5991 3776 6007 3840
rect 6071 3776 6087 3840
rect 6151 3776 6159 3840
rect 5839 2752 6159 3776
rect 5839 2688 5847 2752
rect 5911 2688 5927 2752
rect 5991 2688 6007 2752
rect 6071 2688 6087 2752
rect 6151 2688 6159 2752
rect 5839 2128 6159 2688
rect 7471 45728 7791 46752
rect 7471 45664 7479 45728
rect 7543 45664 7559 45728
rect 7623 45664 7639 45728
rect 7703 45664 7719 45728
rect 7783 45664 7791 45728
rect 7471 44640 7791 45664
rect 7471 44576 7479 44640
rect 7543 44576 7559 44640
rect 7623 44576 7639 44640
rect 7703 44576 7719 44640
rect 7783 44576 7791 44640
rect 7471 43552 7791 44576
rect 7471 43488 7479 43552
rect 7543 43488 7559 43552
rect 7623 43488 7639 43552
rect 7703 43488 7719 43552
rect 7783 43488 7791 43552
rect 7471 42464 7791 43488
rect 7471 42400 7479 42464
rect 7543 42400 7559 42464
rect 7623 42400 7639 42464
rect 7703 42400 7719 42464
rect 7783 42400 7791 42464
rect 7471 41376 7791 42400
rect 7471 41312 7479 41376
rect 7543 41312 7559 41376
rect 7623 41312 7639 41376
rect 7703 41312 7719 41376
rect 7783 41312 7791 41376
rect 7471 40288 7791 41312
rect 7471 40224 7479 40288
rect 7543 40224 7559 40288
rect 7623 40224 7639 40288
rect 7703 40224 7719 40288
rect 7783 40224 7791 40288
rect 7471 39200 7791 40224
rect 7471 39136 7479 39200
rect 7543 39136 7559 39200
rect 7623 39136 7639 39200
rect 7703 39136 7719 39200
rect 7783 39136 7791 39200
rect 7471 38112 7791 39136
rect 7471 38048 7479 38112
rect 7543 38048 7559 38112
rect 7623 38048 7639 38112
rect 7703 38048 7719 38112
rect 7783 38048 7791 38112
rect 7471 37024 7791 38048
rect 7471 36960 7479 37024
rect 7543 36960 7559 37024
rect 7623 36960 7639 37024
rect 7703 36960 7719 37024
rect 7783 36960 7791 37024
rect 7471 35936 7791 36960
rect 7471 35872 7479 35936
rect 7543 35872 7559 35936
rect 7623 35872 7639 35936
rect 7703 35872 7719 35936
rect 7783 35872 7791 35936
rect 7471 34848 7791 35872
rect 7471 34784 7479 34848
rect 7543 34784 7559 34848
rect 7623 34784 7639 34848
rect 7703 34784 7719 34848
rect 7783 34784 7791 34848
rect 7471 33760 7791 34784
rect 7471 33696 7479 33760
rect 7543 33696 7559 33760
rect 7623 33696 7639 33760
rect 7703 33696 7719 33760
rect 7783 33696 7791 33760
rect 7471 32672 7791 33696
rect 7471 32608 7479 32672
rect 7543 32608 7559 32672
rect 7623 32608 7639 32672
rect 7703 32608 7719 32672
rect 7783 32608 7791 32672
rect 7471 31584 7791 32608
rect 7471 31520 7479 31584
rect 7543 31520 7559 31584
rect 7623 31520 7639 31584
rect 7703 31520 7719 31584
rect 7783 31520 7791 31584
rect 7471 30496 7791 31520
rect 7471 30432 7479 30496
rect 7543 30432 7559 30496
rect 7623 30432 7639 30496
rect 7703 30432 7719 30496
rect 7783 30432 7791 30496
rect 7471 29408 7791 30432
rect 7471 29344 7479 29408
rect 7543 29344 7559 29408
rect 7623 29344 7639 29408
rect 7703 29344 7719 29408
rect 7783 29344 7791 29408
rect 7471 28320 7791 29344
rect 7471 28256 7479 28320
rect 7543 28256 7559 28320
rect 7623 28256 7639 28320
rect 7703 28256 7719 28320
rect 7783 28256 7791 28320
rect 7471 27232 7791 28256
rect 7471 27168 7479 27232
rect 7543 27168 7559 27232
rect 7623 27168 7639 27232
rect 7703 27168 7719 27232
rect 7783 27168 7791 27232
rect 7471 26144 7791 27168
rect 7471 26080 7479 26144
rect 7543 26080 7559 26144
rect 7623 26080 7639 26144
rect 7703 26080 7719 26144
rect 7783 26080 7791 26144
rect 7471 25056 7791 26080
rect 7471 24992 7479 25056
rect 7543 24992 7559 25056
rect 7623 24992 7639 25056
rect 7703 24992 7719 25056
rect 7783 24992 7791 25056
rect 7471 23968 7791 24992
rect 7471 23904 7479 23968
rect 7543 23904 7559 23968
rect 7623 23904 7639 23968
rect 7703 23904 7719 23968
rect 7783 23904 7791 23968
rect 7471 22880 7791 23904
rect 7471 22816 7479 22880
rect 7543 22816 7559 22880
rect 7623 22816 7639 22880
rect 7703 22816 7719 22880
rect 7783 22816 7791 22880
rect 7471 21792 7791 22816
rect 7471 21728 7479 21792
rect 7543 21728 7559 21792
rect 7623 21728 7639 21792
rect 7703 21728 7719 21792
rect 7783 21728 7791 21792
rect 7471 20704 7791 21728
rect 7471 20640 7479 20704
rect 7543 20640 7559 20704
rect 7623 20640 7639 20704
rect 7703 20640 7719 20704
rect 7783 20640 7791 20704
rect 7471 19616 7791 20640
rect 7471 19552 7479 19616
rect 7543 19552 7559 19616
rect 7623 19552 7639 19616
rect 7703 19552 7719 19616
rect 7783 19552 7791 19616
rect 7471 18528 7791 19552
rect 7471 18464 7479 18528
rect 7543 18464 7559 18528
rect 7623 18464 7639 18528
rect 7703 18464 7719 18528
rect 7783 18464 7791 18528
rect 7471 17440 7791 18464
rect 7471 17376 7479 17440
rect 7543 17376 7559 17440
rect 7623 17376 7639 17440
rect 7703 17376 7719 17440
rect 7783 17376 7791 17440
rect 7471 16352 7791 17376
rect 7471 16288 7479 16352
rect 7543 16288 7559 16352
rect 7623 16288 7639 16352
rect 7703 16288 7719 16352
rect 7783 16288 7791 16352
rect 7471 15264 7791 16288
rect 7471 15200 7479 15264
rect 7543 15200 7559 15264
rect 7623 15200 7639 15264
rect 7703 15200 7719 15264
rect 7783 15200 7791 15264
rect 7471 14176 7791 15200
rect 7471 14112 7479 14176
rect 7543 14112 7559 14176
rect 7623 14112 7639 14176
rect 7703 14112 7719 14176
rect 7783 14112 7791 14176
rect 7471 13088 7791 14112
rect 7471 13024 7479 13088
rect 7543 13024 7559 13088
rect 7623 13024 7639 13088
rect 7703 13024 7719 13088
rect 7783 13024 7791 13088
rect 7471 12000 7791 13024
rect 7471 11936 7479 12000
rect 7543 11936 7559 12000
rect 7623 11936 7639 12000
rect 7703 11936 7719 12000
rect 7783 11936 7791 12000
rect 7471 10912 7791 11936
rect 7471 10848 7479 10912
rect 7543 10848 7559 10912
rect 7623 10848 7639 10912
rect 7703 10848 7719 10912
rect 7783 10848 7791 10912
rect 7471 9824 7791 10848
rect 7471 9760 7479 9824
rect 7543 9760 7559 9824
rect 7623 9760 7639 9824
rect 7703 9760 7719 9824
rect 7783 9760 7791 9824
rect 7471 8736 7791 9760
rect 7471 8672 7479 8736
rect 7543 8672 7559 8736
rect 7623 8672 7639 8736
rect 7703 8672 7719 8736
rect 7783 8672 7791 8736
rect 7471 7648 7791 8672
rect 7471 7584 7479 7648
rect 7543 7584 7559 7648
rect 7623 7584 7639 7648
rect 7703 7584 7719 7648
rect 7783 7584 7791 7648
rect 7471 6560 7791 7584
rect 7471 6496 7479 6560
rect 7543 6496 7559 6560
rect 7623 6496 7639 6560
rect 7703 6496 7719 6560
rect 7783 6496 7791 6560
rect 7471 5472 7791 6496
rect 7471 5408 7479 5472
rect 7543 5408 7559 5472
rect 7623 5408 7639 5472
rect 7703 5408 7719 5472
rect 7783 5408 7791 5472
rect 7471 4384 7791 5408
rect 7471 4320 7479 4384
rect 7543 4320 7559 4384
rect 7623 4320 7639 4384
rect 7703 4320 7719 4384
rect 7783 4320 7791 4384
rect 7471 3296 7791 4320
rect 7471 3232 7479 3296
rect 7543 3232 7559 3296
rect 7623 3232 7639 3296
rect 7703 3232 7719 3296
rect 7783 3232 7791 3296
rect 7471 2208 7791 3232
rect 7471 2144 7479 2208
rect 7543 2144 7559 2208
rect 7623 2144 7639 2208
rect 7703 2144 7719 2208
rect 7783 2144 7791 2208
rect 7471 2128 7791 2144
rect 9103 77824 9423 77840
rect 9103 77760 9111 77824
rect 9175 77760 9191 77824
rect 9255 77760 9271 77824
rect 9335 77760 9351 77824
rect 9415 77760 9423 77824
rect 9103 76736 9423 77760
rect 9103 76672 9111 76736
rect 9175 76672 9191 76736
rect 9255 76672 9271 76736
rect 9335 76672 9351 76736
rect 9415 76672 9423 76736
rect 9103 75648 9423 76672
rect 9103 75584 9111 75648
rect 9175 75584 9191 75648
rect 9255 75584 9271 75648
rect 9335 75584 9351 75648
rect 9415 75584 9423 75648
rect 9103 74560 9423 75584
rect 9103 74496 9111 74560
rect 9175 74496 9191 74560
rect 9255 74496 9271 74560
rect 9335 74496 9351 74560
rect 9415 74496 9423 74560
rect 9103 73472 9423 74496
rect 9103 73408 9111 73472
rect 9175 73408 9191 73472
rect 9255 73408 9271 73472
rect 9335 73408 9351 73472
rect 9415 73408 9423 73472
rect 9103 72384 9423 73408
rect 9103 72320 9111 72384
rect 9175 72320 9191 72384
rect 9255 72320 9271 72384
rect 9335 72320 9351 72384
rect 9415 72320 9423 72384
rect 9103 71296 9423 72320
rect 9103 71232 9111 71296
rect 9175 71232 9191 71296
rect 9255 71232 9271 71296
rect 9335 71232 9351 71296
rect 9415 71232 9423 71296
rect 9103 70208 9423 71232
rect 9103 70144 9111 70208
rect 9175 70144 9191 70208
rect 9255 70144 9271 70208
rect 9335 70144 9351 70208
rect 9415 70144 9423 70208
rect 9103 69120 9423 70144
rect 9103 69056 9111 69120
rect 9175 69056 9191 69120
rect 9255 69056 9271 69120
rect 9335 69056 9351 69120
rect 9415 69056 9423 69120
rect 9103 68032 9423 69056
rect 9103 67968 9111 68032
rect 9175 67968 9191 68032
rect 9255 67968 9271 68032
rect 9335 67968 9351 68032
rect 9415 67968 9423 68032
rect 9103 66944 9423 67968
rect 9103 66880 9111 66944
rect 9175 66880 9191 66944
rect 9255 66880 9271 66944
rect 9335 66880 9351 66944
rect 9415 66880 9423 66944
rect 9103 65856 9423 66880
rect 9103 65792 9111 65856
rect 9175 65792 9191 65856
rect 9255 65792 9271 65856
rect 9335 65792 9351 65856
rect 9415 65792 9423 65856
rect 9103 64768 9423 65792
rect 9103 64704 9111 64768
rect 9175 64704 9191 64768
rect 9255 64704 9271 64768
rect 9335 64704 9351 64768
rect 9415 64704 9423 64768
rect 9103 63680 9423 64704
rect 9103 63616 9111 63680
rect 9175 63616 9191 63680
rect 9255 63616 9271 63680
rect 9335 63616 9351 63680
rect 9415 63616 9423 63680
rect 9103 62592 9423 63616
rect 9103 62528 9111 62592
rect 9175 62528 9191 62592
rect 9255 62528 9271 62592
rect 9335 62528 9351 62592
rect 9415 62528 9423 62592
rect 9103 61504 9423 62528
rect 9103 61440 9111 61504
rect 9175 61440 9191 61504
rect 9255 61440 9271 61504
rect 9335 61440 9351 61504
rect 9415 61440 9423 61504
rect 9103 60416 9423 61440
rect 9103 60352 9111 60416
rect 9175 60352 9191 60416
rect 9255 60352 9271 60416
rect 9335 60352 9351 60416
rect 9415 60352 9423 60416
rect 9103 59328 9423 60352
rect 9103 59264 9111 59328
rect 9175 59264 9191 59328
rect 9255 59264 9271 59328
rect 9335 59264 9351 59328
rect 9415 59264 9423 59328
rect 9103 58240 9423 59264
rect 9103 58176 9111 58240
rect 9175 58176 9191 58240
rect 9255 58176 9271 58240
rect 9335 58176 9351 58240
rect 9415 58176 9423 58240
rect 9103 57152 9423 58176
rect 9103 57088 9111 57152
rect 9175 57088 9191 57152
rect 9255 57088 9271 57152
rect 9335 57088 9351 57152
rect 9415 57088 9423 57152
rect 9103 56064 9423 57088
rect 9103 56000 9111 56064
rect 9175 56000 9191 56064
rect 9255 56000 9271 56064
rect 9335 56000 9351 56064
rect 9415 56000 9423 56064
rect 9103 54976 9423 56000
rect 9103 54912 9111 54976
rect 9175 54912 9191 54976
rect 9255 54912 9271 54976
rect 9335 54912 9351 54976
rect 9415 54912 9423 54976
rect 9103 53888 9423 54912
rect 9103 53824 9111 53888
rect 9175 53824 9191 53888
rect 9255 53824 9271 53888
rect 9335 53824 9351 53888
rect 9415 53824 9423 53888
rect 9103 52800 9423 53824
rect 9103 52736 9111 52800
rect 9175 52736 9191 52800
rect 9255 52736 9271 52800
rect 9335 52736 9351 52800
rect 9415 52736 9423 52800
rect 9103 51712 9423 52736
rect 9103 51648 9111 51712
rect 9175 51648 9191 51712
rect 9255 51648 9271 51712
rect 9335 51648 9351 51712
rect 9415 51648 9423 51712
rect 9103 50624 9423 51648
rect 9103 50560 9111 50624
rect 9175 50560 9191 50624
rect 9255 50560 9271 50624
rect 9335 50560 9351 50624
rect 9415 50560 9423 50624
rect 9103 49536 9423 50560
rect 9103 49472 9111 49536
rect 9175 49472 9191 49536
rect 9255 49472 9271 49536
rect 9335 49472 9351 49536
rect 9415 49472 9423 49536
rect 9103 48448 9423 49472
rect 9103 48384 9111 48448
rect 9175 48384 9191 48448
rect 9255 48384 9271 48448
rect 9335 48384 9351 48448
rect 9415 48384 9423 48448
rect 9103 47360 9423 48384
rect 9103 47296 9111 47360
rect 9175 47296 9191 47360
rect 9255 47296 9271 47360
rect 9335 47296 9351 47360
rect 9415 47296 9423 47360
rect 9103 46272 9423 47296
rect 9103 46208 9111 46272
rect 9175 46208 9191 46272
rect 9255 46208 9271 46272
rect 9335 46208 9351 46272
rect 9415 46208 9423 46272
rect 9103 45184 9423 46208
rect 9103 45120 9111 45184
rect 9175 45120 9191 45184
rect 9255 45120 9271 45184
rect 9335 45120 9351 45184
rect 9415 45120 9423 45184
rect 9103 44096 9423 45120
rect 9103 44032 9111 44096
rect 9175 44032 9191 44096
rect 9255 44032 9271 44096
rect 9335 44032 9351 44096
rect 9415 44032 9423 44096
rect 9103 43008 9423 44032
rect 9103 42944 9111 43008
rect 9175 42944 9191 43008
rect 9255 42944 9271 43008
rect 9335 42944 9351 43008
rect 9415 42944 9423 43008
rect 9103 41920 9423 42944
rect 9103 41856 9111 41920
rect 9175 41856 9191 41920
rect 9255 41856 9271 41920
rect 9335 41856 9351 41920
rect 9415 41856 9423 41920
rect 9103 40832 9423 41856
rect 9103 40768 9111 40832
rect 9175 40768 9191 40832
rect 9255 40768 9271 40832
rect 9335 40768 9351 40832
rect 9415 40768 9423 40832
rect 9103 39744 9423 40768
rect 9103 39680 9111 39744
rect 9175 39680 9191 39744
rect 9255 39680 9271 39744
rect 9335 39680 9351 39744
rect 9415 39680 9423 39744
rect 9103 38656 9423 39680
rect 9103 38592 9111 38656
rect 9175 38592 9191 38656
rect 9255 38592 9271 38656
rect 9335 38592 9351 38656
rect 9415 38592 9423 38656
rect 9103 37568 9423 38592
rect 9103 37504 9111 37568
rect 9175 37504 9191 37568
rect 9255 37504 9271 37568
rect 9335 37504 9351 37568
rect 9415 37504 9423 37568
rect 9103 36480 9423 37504
rect 9103 36416 9111 36480
rect 9175 36416 9191 36480
rect 9255 36416 9271 36480
rect 9335 36416 9351 36480
rect 9415 36416 9423 36480
rect 9103 35392 9423 36416
rect 9103 35328 9111 35392
rect 9175 35328 9191 35392
rect 9255 35328 9271 35392
rect 9335 35328 9351 35392
rect 9415 35328 9423 35392
rect 9103 34304 9423 35328
rect 9103 34240 9111 34304
rect 9175 34240 9191 34304
rect 9255 34240 9271 34304
rect 9335 34240 9351 34304
rect 9415 34240 9423 34304
rect 9103 33216 9423 34240
rect 9103 33152 9111 33216
rect 9175 33152 9191 33216
rect 9255 33152 9271 33216
rect 9335 33152 9351 33216
rect 9415 33152 9423 33216
rect 9103 32128 9423 33152
rect 9103 32064 9111 32128
rect 9175 32064 9191 32128
rect 9255 32064 9271 32128
rect 9335 32064 9351 32128
rect 9415 32064 9423 32128
rect 9103 31040 9423 32064
rect 9103 30976 9111 31040
rect 9175 30976 9191 31040
rect 9255 30976 9271 31040
rect 9335 30976 9351 31040
rect 9415 30976 9423 31040
rect 9103 29952 9423 30976
rect 9103 29888 9111 29952
rect 9175 29888 9191 29952
rect 9255 29888 9271 29952
rect 9335 29888 9351 29952
rect 9415 29888 9423 29952
rect 9103 28864 9423 29888
rect 9103 28800 9111 28864
rect 9175 28800 9191 28864
rect 9255 28800 9271 28864
rect 9335 28800 9351 28864
rect 9415 28800 9423 28864
rect 9103 27776 9423 28800
rect 9103 27712 9111 27776
rect 9175 27712 9191 27776
rect 9255 27712 9271 27776
rect 9335 27712 9351 27776
rect 9415 27712 9423 27776
rect 9103 26688 9423 27712
rect 9103 26624 9111 26688
rect 9175 26624 9191 26688
rect 9255 26624 9271 26688
rect 9335 26624 9351 26688
rect 9415 26624 9423 26688
rect 9103 25600 9423 26624
rect 9103 25536 9111 25600
rect 9175 25536 9191 25600
rect 9255 25536 9271 25600
rect 9335 25536 9351 25600
rect 9415 25536 9423 25600
rect 9103 24512 9423 25536
rect 9103 24448 9111 24512
rect 9175 24448 9191 24512
rect 9255 24448 9271 24512
rect 9335 24448 9351 24512
rect 9415 24448 9423 24512
rect 9103 23424 9423 24448
rect 9103 23360 9111 23424
rect 9175 23360 9191 23424
rect 9255 23360 9271 23424
rect 9335 23360 9351 23424
rect 9415 23360 9423 23424
rect 9103 22336 9423 23360
rect 9103 22272 9111 22336
rect 9175 22272 9191 22336
rect 9255 22272 9271 22336
rect 9335 22272 9351 22336
rect 9415 22272 9423 22336
rect 9103 21248 9423 22272
rect 9103 21184 9111 21248
rect 9175 21184 9191 21248
rect 9255 21184 9271 21248
rect 9335 21184 9351 21248
rect 9415 21184 9423 21248
rect 9103 20160 9423 21184
rect 9103 20096 9111 20160
rect 9175 20096 9191 20160
rect 9255 20096 9271 20160
rect 9335 20096 9351 20160
rect 9415 20096 9423 20160
rect 9103 19072 9423 20096
rect 9103 19008 9111 19072
rect 9175 19008 9191 19072
rect 9255 19008 9271 19072
rect 9335 19008 9351 19072
rect 9415 19008 9423 19072
rect 9103 17984 9423 19008
rect 9103 17920 9111 17984
rect 9175 17920 9191 17984
rect 9255 17920 9271 17984
rect 9335 17920 9351 17984
rect 9415 17920 9423 17984
rect 9103 16896 9423 17920
rect 9103 16832 9111 16896
rect 9175 16832 9191 16896
rect 9255 16832 9271 16896
rect 9335 16832 9351 16896
rect 9415 16832 9423 16896
rect 9103 15808 9423 16832
rect 9103 15744 9111 15808
rect 9175 15744 9191 15808
rect 9255 15744 9271 15808
rect 9335 15744 9351 15808
rect 9415 15744 9423 15808
rect 9103 14720 9423 15744
rect 9103 14656 9111 14720
rect 9175 14656 9191 14720
rect 9255 14656 9271 14720
rect 9335 14656 9351 14720
rect 9415 14656 9423 14720
rect 9103 13632 9423 14656
rect 9103 13568 9111 13632
rect 9175 13568 9191 13632
rect 9255 13568 9271 13632
rect 9335 13568 9351 13632
rect 9415 13568 9423 13632
rect 9103 12544 9423 13568
rect 9103 12480 9111 12544
rect 9175 12480 9191 12544
rect 9255 12480 9271 12544
rect 9335 12480 9351 12544
rect 9415 12480 9423 12544
rect 9103 11456 9423 12480
rect 9103 11392 9111 11456
rect 9175 11392 9191 11456
rect 9255 11392 9271 11456
rect 9335 11392 9351 11456
rect 9415 11392 9423 11456
rect 9103 10368 9423 11392
rect 9103 10304 9111 10368
rect 9175 10304 9191 10368
rect 9255 10304 9271 10368
rect 9335 10304 9351 10368
rect 9415 10304 9423 10368
rect 9103 9280 9423 10304
rect 9103 9216 9111 9280
rect 9175 9216 9191 9280
rect 9255 9216 9271 9280
rect 9335 9216 9351 9280
rect 9415 9216 9423 9280
rect 9103 8192 9423 9216
rect 9103 8128 9111 8192
rect 9175 8128 9191 8192
rect 9255 8128 9271 8192
rect 9335 8128 9351 8192
rect 9415 8128 9423 8192
rect 9103 7104 9423 8128
rect 9103 7040 9111 7104
rect 9175 7040 9191 7104
rect 9255 7040 9271 7104
rect 9335 7040 9351 7104
rect 9415 7040 9423 7104
rect 9103 6016 9423 7040
rect 9103 5952 9111 6016
rect 9175 5952 9191 6016
rect 9255 5952 9271 6016
rect 9335 5952 9351 6016
rect 9415 5952 9423 6016
rect 9103 4928 9423 5952
rect 9103 4864 9111 4928
rect 9175 4864 9191 4928
rect 9255 4864 9271 4928
rect 9335 4864 9351 4928
rect 9415 4864 9423 4928
rect 9103 3840 9423 4864
rect 9103 3776 9111 3840
rect 9175 3776 9191 3840
rect 9255 3776 9271 3840
rect 9335 3776 9351 3840
rect 9415 3776 9423 3840
rect 9103 2752 9423 3776
rect 9103 2688 9111 2752
rect 9175 2688 9191 2752
rect 9255 2688 9271 2752
rect 9335 2688 9351 2752
rect 9415 2688 9423 2752
rect 9103 2128 9423 2688
use sky130_fd_sc_hd__decap_4  FILLER_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635444444
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input116 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1635444444
transform -1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1635444444
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1635444444
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_18
timestamp 1635444444
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1635444444
transform -1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1635444444
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_30
timestamp 1635444444
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1635444444
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_42
timestamp 1635444444
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1635444444
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1635444444
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1635444444
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1635444444
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1635444444
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1635444444
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1635444444
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1635444444
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1635444444
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1635444444
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1635444444
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_93
timestamp 1635444444
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1635444444
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1635444444
transform 1 0 9660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1635444444
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1635444444
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635444444
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635444444
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_6
timestamp 1635444444
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635444444
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1635444444
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1635444444
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1635444444
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1635444444
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1635444444
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1635444444
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1635444444
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1635444444
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1635444444
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1635444444
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1635444444
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1635444444
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1635444444
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635444444
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_6
timestamp 1635444444
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635444444
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1635444444
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_18
timestamp 1635444444
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_30
timestamp 1635444444
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_42
timestamp 1635444444
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1635444444
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1635444444
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1635444444
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1635444444
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1635444444
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_93
timestamp 1635444444
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1635444444
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1635444444
transform 1 0 9844 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635444444
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_6
timestamp 1635444444
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635444444
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1635444444
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_18
timestamp 1635444444
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1635444444
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1635444444
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1635444444
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1635444444
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1635444444
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1635444444
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1635444444
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1635444444
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1635444444
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1635444444
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp 1635444444
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635444444
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1635444444
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635444444
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_14
timestamp 1635444444
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_21
timestamp 1635444444
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1635444444
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_33
timestamp 1635444444
transform 1 0 4140 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_37
timestamp 1635444444
transform 1 0 4508 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_41
timestamp 1635444444
transform 1 0 4876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1635444444
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1635444444
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1635444444
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1635444444
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1635444444
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1635444444
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1635444444
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1635444444
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635444444
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1635444444
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1635444444
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635444444
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635444444
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _083_
timestamp 1635444444
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1635444444
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _276_
timestamp 1635444444
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1635444444
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1635444444
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_14
timestamp 1635444444
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_21
timestamp 1635444444
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1635444444
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1635444444
transform 1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1635444444
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_32
timestamp 1635444444
transform 1 0 4048 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_33
timestamp 1635444444
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_37
timestamp 1635444444
transform 1 0 4508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1635444444
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _095_
timestamp 1635444444
transform -1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _101_
timestamp 1635444444
transform -1 0 4876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _275_
timestamp 1635444444
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1635444444
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_48
timestamp 1635444444
transform 1 0 5520 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_41
timestamp 1635444444
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _097_
timestamp 1635444444
transform -1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_60
timestamp 1635444444
transform 1 0 6624 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1635444444
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1635444444
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1635444444
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_72
timestamp 1635444444
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1635444444
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1635444444
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1635444444
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1635444444
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_97
timestamp 1635444444
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_93
timestamp 1635444444
transform 1 0 9660 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_99
timestamp 1635444444
transform 1 0 10212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1635444444
transform 1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635444444
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635444444
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1635444444
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635444444
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1635444444
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1635444444
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1635444444
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_37
timestamp 1635444444
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1635444444
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _103_
timestamp 1635444444
transform -1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1635444444
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1635444444
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1635444444
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1635444444
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1635444444
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1635444444
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1635444444
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1635444444
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635444444
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1635444444
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635444444
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1635444444
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1635444444
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1635444444
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1635444444
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1635444444
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1635444444
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1635444444
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1635444444
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1635444444
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1635444444
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1635444444
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1635444444
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635444444
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1635444444
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635444444
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1635444444
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1635444444
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1635444444
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_33
timestamp 1635444444
transform 1 0 4140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1635444444
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _106_
timestamp 1635444444
transform -1 0 4140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_45
timestamp 1635444444
transform 1 0 5244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_57
timestamp 1635444444
transform 1 0 6348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_69
timestamp 1635444444
transform 1 0 7452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1635444444
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1635444444
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1635444444
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1635444444
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635444444
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1635444444
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635444444
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1635444444
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1635444444
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1635444444
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1635444444
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1635444444
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1635444444
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1635444444
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1635444444
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1635444444
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1635444444
transform 1 0 9660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1635444444
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1635444444
transform 1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635444444
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1635444444
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635444444
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1635444444
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1635444444
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1635444444
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1635444444
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1635444444
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1635444444
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1635444444
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1635444444
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1635444444
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1635444444
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1635444444
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 1635444444
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635444444
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1635444444
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_10
timestamp 1635444444
transform 1 0 2024 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635444444
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635444444
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1635444444
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1635444444
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1635444444
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_34
timestamp 1635444444
transform 1 0 4232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1635444444
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_34
timestamp 1635444444
transform 1 0 4232 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1635444444
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _108_
timestamp 1635444444
transform -1 0 4232 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _110_
timestamp 1635444444
transform -1 0 4232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1635444444
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_46
timestamp 1635444444
transform 1 0 5336 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 4784 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1635444444
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_58
timestamp 1635444444
transform 1 0 6440 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1635444444
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1635444444
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_70
timestamp 1635444444
transform 1 0 7544 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1635444444
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1635444444
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1635444444
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1635444444
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_93
timestamp 1635444444
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_99
timestamp 1635444444
transform 1 0 10212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1635444444
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1635444444
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635444444
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635444444
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1635444444
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1635444444
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635444444
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2760 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_18
timestamp 1635444444
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1635444444
transform 1 0 3864 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_34
timestamp 1635444444
transform 1 0 4232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _105_
timestamp 1635444444
transform 1 0 4324 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1635444444
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1635444444
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1635444444
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1635444444
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1635444444
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1635444444
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1635444444
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1635444444
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1635444444
transform 1 0 9844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635444444
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_10
timestamp 1635444444
transform 1 0 2024 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_6
timestamp 1635444444
transform 1 0 1656 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635444444
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2116 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1635444444
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1635444444
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1635444444
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_34
timestamp 1635444444
transform 1 0 4232 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1635444444
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _112_
timestamp 1635444444
transform -1 0 4232 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_46
timestamp 1635444444
transform 1 0 5336 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_58
timestamp 1635444444
transform 1 0 6440 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_70
timestamp 1635444444
transform 1 0 7544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1635444444
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1635444444
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1635444444
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1635444444
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635444444
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1635444444
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635444444
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_18
timestamp 1635444444
transform 1 0 2760 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4_1  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2760 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_17_30
timestamp 1635444444
transform 1 0 3864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_34
timestamp 1635444444
transform 1 0 4232 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _114_
timestamp 1635444444
transform -1 0 4232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_46
timestamp 1635444444
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1635444444
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1635444444
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1635444444
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1635444444
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1635444444
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1635444444
transform 1 0 9660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_99
timestamp 1635444444
transform 1 0 10212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1635444444
transform 1 0 9844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635444444
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_8
timestamp 1635444444
transform 1 0 1840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635444444
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _084_
timestamp 1635444444
transform 1 0 2208 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1635444444
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1635444444
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1635444444
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1635444444
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1635444444
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1635444444
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1635444444
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1635444444
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1635444444
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1635444444
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1635444444
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_97
timestamp 1635444444
transform 1 0 10028 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635444444
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_6
timestamp 1635444444
transform 1 0 1656 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_6
timestamp 1635444444
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635444444
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635444444
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1635444444
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1635444444
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1635444444
transform 1 0 2024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_13
timestamp 1635444444
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_25
timestamp 1635444444
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1635444444
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1635444444
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1635444444
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1635444444
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1635444444
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1635444444
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1635444444
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1635444444
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1635444444
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1635444444
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1635444444
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1635444444
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1635444444
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1635444444
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1635444444
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1635444444
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1635444444
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1635444444
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1635444444
transform 1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1635444444
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_97
timestamp 1635444444
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1635444444
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635444444
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635444444
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_6
timestamp 1635444444
transform 1 0 1656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635444444
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1635444444
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1635444444
transform 1 0 2024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_13
timestamp 1635444444
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_25
timestamp 1635444444
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_37
timestamp 1635444444
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1635444444
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1635444444
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1635444444
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1635444444
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1635444444
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1635444444
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1635444444
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_93
timestamp 1635444444
transform 1 0 9660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635444444
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_9
timestamp 1635444444
transform 1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635444444
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _090_
timestamp 1635444444
transform -1 0 1932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_16
timestamp 1635444444
transform 1 0 2576 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1635444444
transform -1 0 2576 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1635444444
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1635444444
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1635444444
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1635444444
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1635444444
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1635444444
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1635444444
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1635444444
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1635444444
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1635444444
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1635444444
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1635444444
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635444444
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_8
timestamp 1635444444
transform 1 0 1840 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635444444
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _088_
timestamp 1635444444
transform 1 0 1380 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_23_20
timestamp 1635444444
transform 1 0 2944 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_32
timestamp 1635444444
transform 1 0 4048 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_44
timestamp 1635444444
transform 1 0 5152 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1635444444
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1635444444
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1635444444
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1635444444
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1635444444
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_93
timestamp 1635444444
transform 1 0 9660 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635444444
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_6
timestamp 1635444444
transform 1 0 1656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635444444
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1635444444
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1635444444
transform 1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_13
timestamp 1635444444
transform 1 0 2300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1635444444
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1635444444
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1635444444
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1635444444
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1635444444
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1635444444
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1635444444
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1635444444
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1635444444
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1635444444
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1635444444
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_99
timestamp 1635444444
transform 1 0 10212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1635444444
transform 1 0 9844 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635444444
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1635444444
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635444444
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1635444444
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1635444444
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_13
timestamp 1635444444
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_25
timestamp 1635444444
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_37
timestamp 1635444444
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp 1635444444
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1635444444
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1635444444
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1635444444
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1635444444
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1635444444
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1635444444
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_93
timestamp 1635444444
transform 1 0 9660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635444444
transform -1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_12
timestamp 1635444444
transform 1 0 2208 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_6
timestamp 1635444444
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635444444
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635444444
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 1635444444
transform -1 0 2300 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1635444444
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1635444444
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_13
timestamp 1635444444
transform 1 0 2300 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_25
timestamp 1635444444
transform 1 0 3404 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1635444444
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_33
timestamp 1635444444
transform 1 0 4140 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_38
timestamp 1635444444
transform 1 0 4600 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1635444444
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _122_
timestamp 1635444444
transform -1 0 4600 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1635444444
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1635444444
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1635444444
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1635444444
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1635444444
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1635444444
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1635444444
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1635444444
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1635444444
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1635444444
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1635444444
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1635444444
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1635444444
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1635444444
transform 1 0 10212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_101
timestamp 1635444444
transform 1 0 10396 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_93
timestamp 1635444444
transform 1 0 9660 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1635444444
transform 1 0 9844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635444444
transform -1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635444444
transform -1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_6
timestamp 1635444444
transform 1 0 1656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635444444
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp 1635444444
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1635444444
transform -1 0 1656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_13
timestamp 1635444444
transform 1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1635444444
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1635444444
transform 1 0 2668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_29
timestamp 1635444444
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_38
timestamp 1635444444
transform 1 0 4600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1635444444
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _118_
timestamp 1635444444
transform -1 0 4600 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_45
timestamp 1635444444
transform 1 0 5244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _120_
timestamp 1635444444
transform -1 0 5244 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_57
timestamp 1635444444
transform 1 0 6348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_69
timestamp 1635444444
transform 1 0 7452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1635444444
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1635444444
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1635444444
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1635444444
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_99
timestamp 1635444444
transform 1 0 10212 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1635444444
transform 1 0 9844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635444444
transform -1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_6
timestamp 1635444444
transform 1 0 1656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635444444
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 1635444444
transform 1 0 2024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1635444444
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1635444444
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_20
timestamp 1635444444
transform 1 0 2944 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1635444444
transform -1 0 2944 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1635444444
transform 1 0 3312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_27
timestamp 1635444444
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_38
timestamp 1635444444
transform 1 0 4600 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _124_
timestamp 1635444444
transform -1 0 4600 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1635444444
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _126_
timestamp 1635444444
transform -1 0 5244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1635444444
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1635444444
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1635444444
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1635444444
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1635444444
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1635444444
transform 1 0 10396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_93
timestamp 1635444444
transform 1 0 9660 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635444444
transform -1 0 10856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1635444444
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_9
timestamp 1635444444
transform 1 0 1932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635444444
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113_
timestamp 1635444444
transform -1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp 1635444444
transform 1 0 3128 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 3128 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1635444444
transform 1 0 4048 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1635444444
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1635444444
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1635444444
transform 1 0 5152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1635444444
transform 1 0 6256 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1635444444
transform 1 0 7360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1635444444
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1635444444
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1635444444
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1635444444
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 1635444444
transform 1 0 10212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1635444444
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635444444
transform -1 0 10856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1635444444
transform 1 0 1380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1635444444
transform 1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635444444
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 1932 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_31_22
timestamp 1635444444
transform 1 0 3128 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _197_
timestamp 1635444444
transform -1 0 3128 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_31_31
timestamp 1635444444
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _196_
timestamp 1635444444
transform -1 0 3956 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_31_43
timestamp 1635444444
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1635444444
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1635444444
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1635444444
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1635444444
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1635444444
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_101
timestamp 1635444444
transform 1 0 10396 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_93
timestamp 1635444444
transform 1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635444444
transform -1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1635444444
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1635444444
transform 1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635444444
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1635444444
transform -1 0 1932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_18
timestamp 1635444444
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _194_
timestamp 1635444444
transform -1 0 2760 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1635444444
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1635444444
transform 1 0 4048 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1635444444
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1635444444
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1635444444
transform 1 0 5152 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1635444444
transform 1 0 6256 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1635444444
transform 1 0 7360 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1635444444
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1635444444
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1635444444
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1635444444
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1635444444
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1635444444
transform 1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635444444
transform -1 0 10856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_6
timestamp 1635444444
transform 1 0 1656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_6
timestamp 1635444444
transform 1 0 1656 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635444444
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635444444
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1635444444
transform -1 0 2300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1635444444
transform -1 0 1656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1635444444
transform 1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1635444444
transform -1 0 1656 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_13
timestamp 1635444444
transform 1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_20
timestamp 1635444444
transform 1 0 2944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_13
timestamp 1635444444
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_17
timestamp 1635444444
transform 1 0 2668 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1635444444
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 1635444444
transform 1 0 2668 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _193_
timestamp 1635444444
transform -1 0 3128 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1635444444
transform 1 0 3312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1635444444
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp 1635444444
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_35
timestamp 1635444444
transform 1 0 4324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1635444444
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _117_
timestamp 1635444444
transform 1 0 4416 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1635444444
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1635444444
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_46
timestamp 1635444444
transform 1 0 5336 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1635444444
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1635444444
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_58
timestamp 1635444444
transform 1 0 6440 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1635444444
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1635444444
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_70
timestamp 1635444444
transform 1 0 7544 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1635444444
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1635444444
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1635444444
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1635444444
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_101
timestamp 1635444444
transform 1 0 10396 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_93
timestamp 1635444444
transform 1 0 9660 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1635444444
transform 1 0 9660 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1635444444
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1635444444
transform 1 0 9844 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635444444
transform -1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635444444
transform -1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_6
timestamp 1635444444
transform 1 0 1656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635444444
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1635444444
transform 1 0 2024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1635444444
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_13
timestamp 1635444444
transform 1 0 2300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_20
timestamp 1635444444
transform 1 0 2944 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1635444444
transform 1 0 2668 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1635444444
transform -1 0 3588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1635444444
transform 1 0 3588 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_31
timestamp 1635444444
transform 1 0 3956 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_35
timestamp 1635444444
transform 1 0 4324 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _129_
timestamp 1635444444
transform -1 0 4324 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_42
timestamp 1635444444
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _131_
timestamp 1635444444
transform -1 0 4968 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1635444444
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1635444444
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1635444444
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1635444444
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1635444444
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_101
timestamp 1635444444
transform 1 0 10396 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_93
timestamp 1635444444
transform 1 0 9660 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635444444
transform -1 0 10856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_6
timestamp 1635444444
transform 1 0 1656 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635444444
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _127_
timestamp 1635444444
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1635444444
transform -1 0 2300 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1635444444
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_17
timestamp 1635444444
transform 1 0 2668 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_22
timestamp 1635444444
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 3128 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_29
timestamp 1635444444
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_35
timestamp 1635444444
transform 1 0 4324 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1635444444
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _133_
timestamp 1635444444
transform -1 0 4324 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_47
timestamp 1635444444
transform 1 0 5428 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_59
timestamp 1635444444
transform 1 0 6532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_71
timestamp 1635444444
transform 1 0 7636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1635444444
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1635444444
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1635444444
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1635444444
transform 1 0 9660 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1635444444
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1635444444
transform 1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635444444
transform -1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_6
timestamp 1635444444
transform 1 0 1656 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635444444
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _130_
timestamp 1635444444
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _200_
timestamp 1635444444
transform 1 0 2024 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_37_15
timestamp 1635444444
transform 1 0 2484 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_24
timestamp 1635444444
transform 1 0 3312 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _201_
timestamp 1635444444
transform -1 0 3312 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_37_32
timestamp 1635444444
transform 1 0 4048 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1635444444
transform 1 0 4232 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_37_44
timestamp 1635444444
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1635444444
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1635444444
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1635444444
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1635444444
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_101
timestamp 1635444444
transform 1 0 10396 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_93
timestamp 1635444444
transform 1 0 9660 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635444444
transform -1 0 10856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_6
timestamp 1635444444
transform 1 0 1656 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635444444
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _132_
timestamp 1635444444
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _202_
timestamp 1635444444
transform -1 0 2484 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_38_15
timestamp 1635444444
transform 1 0 2484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 1635444444
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1635444444
transform 1 0 2852 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1635444444
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1635444444
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_35
timestamp 1635444444
transform 1 0 4324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1635444444
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _135_
timestamp 1635444444
transform -1 0 4324 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_42
timestamp 1635444444
transform 1 0 4968 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _137_
timestamp 1635444444
transform -1 0 4968 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_54
timestamp 1635444444
transform 1 0 6072 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_66
timestamp 1635444444
transform 1 0 7176 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_78
timestamp 1635444444
transform 1 0 8280 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_85
timestamp 1635444444
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1635444444
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1635444444
transform 1 0 9660 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_99
timestamp 1635444444
transform 1 0 10212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1635444444
transform 1 0 9844 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635444444
transform -1 0 10856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1635444444
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_6
timestamp 1635444444
transform 1 0 1656 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635444444
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635444444
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _134_
timestamp 1635444444
transform -1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1635444444
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _203_
timestamp 1635444444
transform 1 0 1932 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1635444444
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_23
timestamp 1635444444
transform 1 0 3220 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_13
timestamp 1635444444
transform 1 0 2300 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1635444444
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _204_
timestamp 1635444444
transform -1 0 3220 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1635444444
transform 1 0 2668 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_30
timestamp 1635444444
transform 1 0 3864 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1635444444
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_37
timestamp 1635444444
transform 1 0 4508 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1635444444
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1635444444
transform 1 0 4140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1635444444
transform 1 0 3588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_42
timestamp 1635444444
transform 1 0 4968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_49
timestamp 1635444444
transform 1 0 5612 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1635444444
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1635444444
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_61
timestamp 1635444444
transform 1 0 6716 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1635444444
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1635444444
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_73
timestamp 1635444444
transform 1 0 7820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1635444444
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 1635444444
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1635444444
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1635444444
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_101
timestamp 1635444444
transform 1 0 10396 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_93
timestamp 1635444444
transform 1 0 9660 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1635444444
transform 1 0 9660 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1635444444
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1635444444
transform 1 0 9844 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635444444
transform -1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635444444
transform -1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_6
timestamp 1635444444
transform 1 0 1656 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635444444
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1635444444
transform -1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_18
timestamp 1635444444
transform 1 0 2760 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_22
timestamp 1635444444
transform 1 0 3128 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1635444444
transform 1 0 3220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_26
timestamp 1635444444
transform 1 0 3496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_30
timestamp 1635444444
transform 1 0 3864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_37
timestamp 1635444444
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1635444444
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1635444444
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1635444444
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1635444444
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1635444444
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1635444444
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_101
timestamp 1635444444
transform 1 0 10396 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_93
timestamp 1635444444
transform 1 0 9660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635444444
transform -1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_6
timestamp 1635444444
transform 1 0 1656 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635444444
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1635444444
transform -1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1635444444
transform 1 0 2024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_13
timestamp 1635444444
transform 1 0 2300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1635444444
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1635444444
transform 1 0 2668 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1635444444
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1635444444
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1635444444
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1635444444
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1635444444
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1635444444
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1635444444
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1635444444
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1635444444
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 1635444444
transform 1 0 9660 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1635444444
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1635444444
transform 1 0 9844 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635444444
transform -1 0 10856 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_6
timestamp 1635444444
transform 1 0 1656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635444444
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1635444444
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1635444444
transform 1 0 2024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_13
timestamp 1635444444
transform 1 0 2300 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_25
timestamp 1635444444
transform 1 0 3404 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_37
timestamp 1635444444
transform 1 0 4508 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_49
timestamp 1635444444
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1635444444
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1635444444
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1635444444
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1635444444
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1635444444
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_101
timestamp 1635444444
transform 1 0 10396 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1635444444
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635444444
transform -1 0 10856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_6
timestamp 1635444444
transform 1 0 1656 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635444444
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp 1635444444
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1635444444
transform -1 0 2300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_13
timestamp 1635444444
transform 1 0 2300 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_17
timestamp 1635444444
transform 1 0 2668 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1635444444
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _229_
timestamp 1635444444
transform -1 0 3312 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_32
timestamp 1635444444
transform 1 0 4048 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1635444444
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _140_
timestamp 1635444444
transform -1 0 4048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _142_
timestamp 1635444444
transform -1 0 4692 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_39
timestamp 1635444444
transform 1 0 4692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_51
timestamp 1635444444
transform 1 0 5796 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_63
timestamp 1635444444
transform 1 0 6900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_75
timestamp 1635444444
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1635444444
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_85
timestamp 1635444444
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1635444444
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_93
timestamp 1635444444
transform 1 0 9660 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_99
timestamp 1635444444
transform 1 0 10212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1635444444
transform 1 0 9844 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635444444
transform -1 0 10856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_6
timestamp 1635444444
transform 1 0 1656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635444444
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1635444444
transform -1 0 1656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1635444444
transform 1 0 2024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_13
timestamp 1635444444
transform 1 0 2300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_20
timestamp 1635444444
transform 1 0 2944 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1635444444
transform 1 0 2668 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_26
timestamp 1635444444
transform 1 0 3496 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_30
timestamp 1635444444
transform 1 0 3864 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _144_
timestamp 1635444444
transform -1 0 3864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_42
timestamp 1635444444
transform 1 0 4968 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1635444444
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1635444444
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1635444444
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1635444444
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1635444444
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_101
timestamp 1635444444
transform 1 0 10396 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_93
timestamp 1635444444
transform 1 0 9660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635444444
transform -1 0 10856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_6
timestamp 1635444444
transform 1 0 1656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1635444444
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_7
timestamp 1635444444
transform 1 0 1748 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635444444
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1635444444
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1635444444
transform -1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _206_
timestamp 1635444444
transform 1 0 1840 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1635444444
transform 1 0 2024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_13
timestamp 1635444444
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_17
timestamp 1635444444
transform 1 0 2668 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_22
timestamp 1635444444
transform 1 0 3128 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_13
timestamp 1635444444
transform 1 0 2300 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_22
timestamp 1635444444
transform 1 0 3128 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _205_
timestamp 1635444444
transform -1 0 3128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _207_
timestamp 1635444444
transform -1 0 3128 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1635444444
transform 1 0 4048 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_30
timestamp 1635444444
transform 1 0 3864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1635444444
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _139_
timestamp 1635444444
transform 1 0 3956 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _146_
timestamp 1635444444
transform -1 0 4048 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1635444444
transform 1 0 5152 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_41
timestamp 1635444444
transform 1 0 4876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_56
timestamp 1635444444
transform 1 0 6256 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1635444444
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1635444444
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1635444444
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_68
timestamp 1635444444
transform 1 0 7360 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1635444444
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1635444444
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1635444444
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1635444444
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1635444444
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_93
timestamp 1635444444
transform 1 0 9660 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1635444444
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_101
timestamp 1635444444
transform 1 0 10396 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_93
timestamp 1635444444
transform 1 0 9660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1635444444
transform 1 0 9844 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635444444
transform -1 0 10856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1635444444
transform -1 0 10856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1635444444
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_7
timestamp 1635444444
transform 1 0 1748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1635444444
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _208_
timestamp 1635444444
transform -1 0 2300 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_48_13
timestamp 1635444444
transform 1 0 2300 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_22
timestamp 1635444444
transform 1 0 3128 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _209_
timestamp 1635444444
transform -1 0 3128 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1635444444
transform 1 0 4048 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1635444444
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _148_
timestamp 1635444444
transform -1 0 4048 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1635444444
transform 1 0 5152 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_56
timestamp 1635444444
transform 1 0 6256 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_68
timestamp 1635444444
transform 1 0 7360 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1635444444
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1635444444
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1635444444
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1635444444
transform 1 0 9660 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_99
timestamp 1635444444
transform 1 0 10212 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1635444444
transform 1 0 9844 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1635444444
transform -1 0 10856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1635444444
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_7
timestamp 1635444444
transform 1 0 1748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1635444444
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _210_
timestamp 1635444444
transform -1 0 2300 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_49_13
timestamp 1635444444
transform 1 0 2300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_20
timestamp 1635444444
transform 1 0 2944 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1635444444
transform 1 0 2668 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1635444444
transform 1 0 3312 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1635444444
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1635444444
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1635444444
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1635444444
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1635444444
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1635444444
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1635444444
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1635444444
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_101
timestamp 1635444444
transform 1 0 10396 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_93
timestamp 1635444444
transform 1 0 9660 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1635444444
transform -1 0 10856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_10
timestamp 1635444444
transform 1 0 2024 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1635444444
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1635444444
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _149_
timestamp 1635444444
transform -1 0 2024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_17
timestamp 1635444444
transform 1 0 2668 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1635444444
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1635444444
transform 1 0 3036 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1635444444
transform 1 0 2392 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1635444444
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1635444444
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1635444444
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1635444444
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1635444444
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1635444444
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1635444444
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1635444444
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1635444444
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_93
timestamp 1635444444
transform 1 0 9660 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_99
timestamp 1635444444
transform 1 0 10212 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1635444444
transform 1 0 9844 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1635444444
transform -1 0 10856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_3
timestamp 1635444444
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_9
timestamp 1635444444
transform 1 0 1932 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1635444444
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152_
timestamp 1635444444
transform -1 0 1932 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_16
timestamp 1635444444
transform 1 0 2576 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1635444444
transform -1 0 2576 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_28
timestamp 1635444444
transform 1 0 3680 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_40
timestamp 1635444444
transform 1 0 4784 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1635444444
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1635444444
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1635444444
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1635444444
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1635444444
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_101
timestamp 1635444444
transform 1 0 10396 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_93
timestamp 1635444444
transform 1 0 9660 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1635444444
transform -1 0 10856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_3
timestamp 1635444444
transform 1 0 1380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_9
timestamp 1635444444
transform 1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_3
timestamp 1635444444
transform 1 0 1380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_9
timestamp 1635444444
transform 1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1635444444
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1635444444
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1635444444
transform -1 0 1932 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 1635444444
transform -1 0 1932 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_16
timestamp 1635444444
transform 1 0 2576 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_23
timestamp 1635444444
transform 1 0 3220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_16
timestamp 1635444444
transform 1 0 2576 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp 1635444444
transform 1 0 2300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1635444444
transform 1 0 2300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1635444444
transform 1 0 2944 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1635444444
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_32
timestamp 1635444444
transform 1 0 4048 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_28
timestamp 1635444444
transform 1 0 3680 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1635444444
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _151_
timestamp 1635444444
transform -1 0 4692 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _153_
timestamp 1635444444
transform -1 0 4692 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1635444444
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_39
timestamp 1635444444
transform 1 0 4692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_51
timestamp 1635444444
transform 1 0 5796 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1635444444
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1635444444
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_63
timestamp 1635444444
transform 1 0 6900 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1635444444
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1635444444
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1635444444
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_75
timestamp 1635444444
transform 1 0 8004 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1635444444
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1635444444
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1635444444
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1635444444
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1635444444
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 1635444444
transform 1 0 9660 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1635444444
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_101
timestamp 1635444444
transform 1 0 10396 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_93
timestamp 1635444444
transform 1 0 9660 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1635444444
transform 1 0 9844 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1635444444
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1635444444
transform -1 0 10856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_11
timestamp 1635444444
transform 1 0 2116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1635444444
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_7
timestamp 1635444444
transform 1 0 1748 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1635444444
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1635444444
transform -1 0 2116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_18
timestamp 1635444444
transform 1 0 2760 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1635444444
transform 1 0 2484 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1635444444
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_29
timestamp 1635444444
transform 1 0 3772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_35
timestamp 1635444444
transform 1 0 4324 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1635444444
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _155_
timestamp 1635444444
transform -1 0 4692 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_39
timestamp 1635444444
transform 1 0 4692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_51
timestamp 1635444444
transform 1 0 5796 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_63
timestamp 1635444444
transform 1 0 6900 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_75
timestamp 1635444444
transform 1 0 8004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1635444444
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1635444444
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1635444444
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_93
timestamp 1635444444
transform 1 0 9660 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_99
timestamp 1635444444
transform 1 0 10212 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1635444444
transform 1 0 9844 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1635444444
transform -1 0 10856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_6
timestamp 1635444444
transform 1 0 1656 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1635444444
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _213_
timestamp 1635444444
transform -1 0 2668 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1635444444
transform -1 0 1656 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_17
timestamp 1635444444
transform 1 0 2668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_25
timestamp 1635444444
transform 1 0 3404 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _211_
timestamp 1635444444
transform 1 0 3036 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_33
timestamp 1635444444
transform 1 0 4140 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _150_
timestamp 1635444444
transform 1 0 4324 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1635444444
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1635444444
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1635444444
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1635444444
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1635444444
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1635444444
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_101
timestamp 1635444444
transform 1 0 10396 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_93
timestamp 1635444444
transform 1 0 9660 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1635444444
transform -1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_11
timestamp 1635444444
transform 1 0 2116 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_7
timestamp 1635444444
transform 1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1635444444
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _212_
timestamp 1635444444
transform -1 0 2668 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1635444444
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_17
timestamp 1635444444
transform 1 0 2668 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1635444444
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1635444444
transform 1 0 3036 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_29
timestamp 1635444444
transform 1 0 3772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_38
timestamp 1635444444
transform 1 0 4600 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1635444444
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _157_
timestamp 1635444444
transform -1 0 4600 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_50
timestamp 1635444444
transform 1 0 5704 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_62
timestamp 1635444444
transform 1 0 6808 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_74
timestamp 1635444444
transform 1 0 7912 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1635444444
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1635444444
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1635444444
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_93
timestamp 1635444444
transform 1 0 9660 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_99
timestamp 1635444444
transform 1 0 10212 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1635444444
transform 1 0 9844 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1635444444
transform -1 0 10856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_3
timestamp 1635444444
transform 1 0 1380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_8
timestamp 1635444444
transform 1 0 1840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1635444444
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 1840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _214_
timestamp 1635444444
transform -1 0 2668 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_57_17
timestamp 1635444444
transform 1 0 2668 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _215_
timestamp 1635444444
transform -1 0 3496 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_57_26
timestamp 1635444444
transform 1 0 3496 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_34
timestamp 1635444444
transform 1 0 4232 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_38
timestamp 1635444444
transform 1 0 4600 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _159_
timestamp 1635444444
transform -1 0 4600 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_50
timestamp 1635444444
transform 1 0 5704 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1635444444
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1635444444
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1635444444
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1635444444
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_101
timestamp 1635444444
transform 1 0 10396 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_93
timestamp 1635444444
transform 1 0 9660 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1635444444
transform -1 0 10856 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_11
timestamp 1635444444
transform 1 0 2116 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_7
timestamp 1635444444
transform 1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1635444444
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _216_
timestamp 1635444444
transform -1 0 2668 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1635444444
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_17
timestamp 1635444444
transform 1 0 2668 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1635444444
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1635444444
transform 1 0 3036 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1635444444
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1635444444
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1635444444
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1635444444
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1635444444
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1635444444
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1635444444
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1635444444
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1635444444
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1635444444
transform 1 0 9660 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_99
timestamp 1635444444
transform 1 0 10212 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1635444444
transform 1 0 9844 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1635444444
transform -1 0 10856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_11
timestamp 1635444444
transform 1 0 2116 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_7
timestamp 1635444444
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_7
timestamp 1635444444
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1635444444
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1635444444
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _173_
timestamp 1635444444
transform -1 0 2576 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1635444444
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1635444444
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_16
timestamp 1635444444
transform 1 0 2576 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_24
timestamp 1635444444
transform 1 0 3312 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 1635444444
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _175_
timestamp 1635444444
transform 1 0 2944 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_36
timestamp 1635444444
transform 1 0 4416 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1635444444
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_29
timestamp 1635444444
transform 1 0 3772 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_33
timestamp 1635444444
transform 1 0 4140 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1635444444
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _161_
timestamp 1635444444
transform 1 0 4232 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_59_48
timestamp 1635444444
transform 1 0 5520 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1635444444
transform 1 0 5152 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1635444444
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_56
timestamp 1635444444
transform 1 0 6256 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1635444444
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1635444444
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_68
timestamp 1635444444
transform 1 0 7360 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1635444444
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1635444444
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_85
timestamp 1635444444
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1635444444
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_101
timestamp 1635444444
transform 1 0 10396 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_93
timestamp 1635444444
transform 1 0 9660 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_93
timestamp 1635444444
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_99
timestamp 1635444444
transform 1 0 10212 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1635444444
transform 1 0 9844 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1635444444
transform -1 0 10856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1635444444
transform -1 0 10856 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1635444444
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1635444444
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1635444444
transform -1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1635444444
transform 1 0 2116 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_15
timestamp 1635444444
transform 1 0 2484 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_23
timestamp 1635444444
transform 1 0 3220 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _217_
timestamp 1635444444
transform -1 0 3220 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_35
timestamp 1635444444
transform 1 0 4324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_47
timestamp 1635444444
transform 1 0 5428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1635444444
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1635444444
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1635444444
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1635444444
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1635444444
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_101
timestamp 1635444444
transform 1 0 10396 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_93
timestamp 1635444444
transform 1 0 9660 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1635444444
transform -1 0 10856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_7
timestamp 1635444444
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1635444444
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1635444444
transform -1 0 2392 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1635444444
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_14
timestamp 1635444444
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1635444444
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_29
timestamp 1635444444
transform 1 0 3772 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_36
timestamp 1635444444
transform 1 0 4416 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1635444444
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _162_
timestamp 1635444444
transform -1 0 4416 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_48
timestamp 1635444444
transform 1 0 5520 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_60
timestamp 1635444444
transform 1 0 6624 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_72
timestamp 1635444444
transform 1 0 7728 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_85
timestamp 1635444444
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1635444444
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_93
timestamp 1635444444
transform 1 0 9660 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_99
timestamp 1635444444
transform 1 0 10212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1635444444
transform 1 0 9844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1635444444
transform -1 0 10856 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_7
timestamp 1635444444
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1635444444
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1635444444
transform -1 0 2392 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1635444444
transform -1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_14
timestamp 1635444444
transform 1 0 2392 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_21
timestamp 1635444444
transform 1 0 3036 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1635444444
transform 1 0 2760 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_36
timestamp 1635444444
transform 1 0 4416 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _164_
timestamp 1635444444
transform -1 0 4416 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_48
timestamp 1635444444
transform 1 0 5520 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1635444444
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1635444444
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1635444444
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1635444444
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_101
timestamp 1635444444
transform 1 0 10396 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_93
timestamp 1635444444
transform 1 0 9660 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1635444444
transform -1 0 10856 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_7
timestamp 1635444444
transform 1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1635444444
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1635444444
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1635444444
transform 1 0 2116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1635444444
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_22
timestamp 1635444444
transform 1 0 3128 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1635444444
transform -1 0 3128 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1635444444
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1635444444
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1635444444
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1635444444
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1635444444
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1635444444
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1635444444
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1635444444
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1635444444
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_93
timestamp 1635444444
transform 1 0 9660 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_99
timestamp 1635444444
transform 1 0 10212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1635444444
transform 1 0 9844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1635444444
transform -1 0 10856 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_65_11
timestamp 1635444444
transform 1 0 2116 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_7
timestamp 1635444444
transform 1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1635444444
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _218_
timestamp 1635444444
transform 1 0 2208 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1635444444
transform -1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_17
timestamp 1635444444
transform 1 0 2668 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_25
timestamp 1635444444
transform 1 0 3404 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1635444444
transform 1 0 3036 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_36
timestamp 1635444444
transform 1 0 4416 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _166_
timestamp 1635444444
transform -1 0 4416 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_48
timestamp 1635444444
transform 1 0 5520 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1635444444
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1635444444
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1635444444
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1635444444
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_101
timestamp 1635444444
transform 1 0 10396 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_93
timestamp 1635444444
transform 1 0 9660 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1635444444
transform -1 0 10856 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_7
timestamp 1635444444
transform 1 0 1748 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_7
timestamp 1635444444
transform 1 0 1748 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1635444444
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1635444444
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1635444444
transform -1 0 1748 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1635444444
transform -1 0 1748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_18
timestamp 1635444444
transform 1 0 2760 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_18
timestamp 1635444444
transform 1 0 2760 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _219_
timestamp 1635444444
transform -1 0 2760 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _220_
timestamp 1635444444
transform -1 0 2760 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_66_26
timestamp 1635444444
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_29
timestamp 1635444444
transform 1 0 3772 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_33
timestamp 1635444444
transform 1 0 4140 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_37
timestamp 1635444444
transform 1 0 4508 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_30
timestamp 1635444444
transform 1 0 3864 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_37
timestamp 1635444444
transform 1 0 4508 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1635444444
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _168_
timestamp 1635444444
transform -1 0 4508 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _170_
timestamp 1635444444
transform -1 0 4508 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_49
timestamp 1635444444
transform 1 0 5612 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_49
timestamp 1635444444
transform 1 0 5612 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_61
timestamp 1635444444
transform 1 0 6716 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1635444444
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1635444444
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1635444444
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_73
timestamp 1635444444
transform 1 0 7820 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1635444444
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_81
timestamp 1635444444
transform 1 0 8556 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_85
timestamp 1635444444
transform 1 0 8924 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1635444444
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1635444444
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_93
timestamp 1635444444
transform 1 0 9660 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_99
timestamp 1635444444
transform 1 0 10212 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_101
timestamp 1635444444
transform 1 0 10396 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_93
timestamp 1635444444
transform 1 0 9660 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1635444444
transform 1 0 9844 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1635444444
transform -1 0 10856 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1635444444
transform -1 0 10856 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_7
timestamp 1635444444
transform 1 0 1748 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1635444444
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1635444444
transform -1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_18
timestamp 1635444444
transform 1 0 2760 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _221_
timestamp 1635444444
transform -1 0 2760 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_68_26
timestamp 1635444444
transform 1 0 3496 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1635444444
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1635444444
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1635444444
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1635444444
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1635444444
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1635444444
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1635444444
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_85
timestamp 1635444444
transform 1 0 8924 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1635444444
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_93
timestamp 1635444444
transform 1 0 9660 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_99
timestamp 1635444444
transform 1 0 10212 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1635444444
transform 1 0 9844 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1635444444
transform -1 0 10856 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_7
timestamp 1635444444
transform 1 0 1748 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1635444444
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1635444444
transform -1 0 1748 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_18
timestamp 1635444444
transform 1 0 2760 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _222_
timestamp 1635444444
transform -1 0 2760 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_69_30
timestamp 1635444444
transform 1 0 3864 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_42
timestamp 1635444444
transform 1 0 4968 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_54
timestamp 1635444444
transform 1 0 6072 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1635444444
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1635444444
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1635444444
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1635444444
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_101
timestamp 1635444444
transform 1 0 10396 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_93
timestamp 1635444444
transform 1 0 9660 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1635444444
transform -1 0 10856 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_7
timestamp 1635444444
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1635444444
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1635444444
transform -1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 1635444444
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1635444444
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1635444444
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1635444444
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1635444444
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1635444444
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1635444444
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1635444444
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1635444444
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1635444444
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1635444444
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_97
timestamp 1635444444
transform 1 0 10028 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1635444444
transform -1 0 10856 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_7
timestamp 1635444444
transform 1 0 1748 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1635444444
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1635444444
transform -1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_19
timestamp 1635444444
transform 1 0 2852 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_31
timestamp 1635444444
transform 1 0 3956 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _172_
timestamp 1635444444
transform -1 0 4784 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_40
timestamp 1635444444
transform 1 0 4784 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_52
timestamp 1635444444
transform 1 0 5888 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1635444444
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1635444444
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1635444444
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1635444444
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_93
timestamp 1635444444
transform 1 0 9660 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_99
timestamp 1635444444
transform 1 0 10212 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1635444444
transform 1 0 9844 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1635444444
transform -1 0 10856 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_7
timestamp 1635444444
transform 1 0 1748 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_7
timestamp 1635444444
transform 1 0 1748 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1635444444
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1635444444
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1635444444
transform -1 0 1748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1635444444
transform -1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_19
timestamp 1635444444
transform 1 0 2852 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_19
timestamp 1635444444
transform 1 0 2852 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1635444444
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1635444444
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_31
timestamp 1635444444
transform 1 0 3956 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1635444444
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _174_
timestamp 1635444444
transform -1 0 4784 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1635444444
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_40
timestamp 1635444444
transform 1 0 4784 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1635444444
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_52
timestamp 1635444444
transform 1 0 5888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1635444444
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1635444444
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1635444444
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1635444444
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1635444444
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1635444444
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1635444444
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1635444444
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1635444444
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_97
timestamp 1635444444
transform 1 0 10028 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_93
timestamp 1635444444
transform 1 0 9660 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_99
timestamp 1635444444
transform 1 0 10212 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1635444444
transform 1 0 9844 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1635444444
transform -1 0 10856 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1635444444
transform -1 0 10856 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_7
timestamp 1635444444
transform 1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1635444444
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1635444444
transform -1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1635444444
transform -1 0 2484 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1635444444
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1635444444
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_29
timestamp 1635444444
transform 1 0 3772 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1635444444
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _176_
timestamp 1635444444
transform -1 0 4784 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_40
timestamp 1635444444
transform 1 0 4784 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_52
timestamp 1635444444
transform 1 0 5888 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_64
timestamp 1635444444
transform 1 0 6992 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_76
timestamp 1635444444
transform 1 0 8096 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1635444444
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1635444444
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_97
timestamp 1635444444
transform 1 0 10028 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1635444444
transform -1 0 10856 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_10
timestamp 1635444444
transform 1 0 2024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1635444444
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2024 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_75_18
timestamp 1635444444
transform 1 0 2760 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1635444444
transform -1 0 2760 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_30
timestamp 1635444444
transform 1 0 3864 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_42
timestamp 1635444444
transform 1 0 4968 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_54
timestamp 1635444444
transform 1 0 6072 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1635444444
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1635444444
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1635444444
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1635444444
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_93
timestamp 1635444444
transform 1 0 9660 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_99
timestamp 1635444444
transform 1 0 10212 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1635444444
transform 1 0 9844 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1635444444
transform -1 0 10856 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_10
timestamp 1635444444
transform 1 0 2024 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1635444444
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _232_
timestamp 1635444444
transform -1 0 2024 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_76_18
timestamp 1635444444
transform 1 0 2760 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1635444444
transform 1 0 2392 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_26
timestamp 1635444444
transform 1 0 3496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_33
timestamp 1635444444
transform 1 0 4140 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1635444444
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1635444444
transform 1 0 3772 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_45
timestamp 1635444444
transform 1 0 5244 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_57
timestamp 1635444444
transform 1 0 6348 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_69
timestamp 1635444444
transform 1 0 7452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_81
timestamp 1635444444
transform 1 0 8556 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1635444444
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1635444444
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_97
timestamp 1635444444
transform 1 0 10028 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1635444444
transform -1 0 10856 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_10
timestamp 1635444444
transform 1 0 2024 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1635444444
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _234_
timestamp 1635444444
transform -1 0 2024 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_77_21
timestamp 1635444444
transform 1 0 3036 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _236_
timestamp 1635444444
transform -1 0 3036 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_77_33
timestamp 1635444444
transform 1 0 4140 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_45
timestamp 1635444444
transform 1 0 5244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1635444444
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1635444444
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1635444444
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1635444444
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1635444444
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_93
timestamp 1635444444
transform 1 0 9660 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_99
timestamp 1635444444
transform 1 0 10212 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1635444444
transform 1 0 9936 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1635444444
transform -1 0 10856 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_10
timestamp 1635444444
transform 1 0 2024 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1635444444
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _235_
timestamp 1635444444
transform -1 0 2024 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_78_18
timestamp 1635444444
transform 1 0 2760 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1635444444
transform -1 0 2760 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_26
timestamp 1635444444
transform 1 0 3496 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1635444444
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1635444444
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1635444444
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1635444444
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1635444444
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1635444444
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1635444444
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1635444444
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1635444444
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_97
timestamp 1635444444
transform 1 0 10028 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1635444444
transform -1 0 10856 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1635444444
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_7
timestamp 1635444444
transform 1 0 1748 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_7
timestamp 1635444444
transform 1 0 1748 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1635444444
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1635444444
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _231_
timestamp 1635444444
transform -1 0 2760 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1635444444
transform -1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_18
timestamp 1635444444
transform 1 0 2760 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_13
timestamp 1635444444
transform 1 0 2300 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1635444444
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _228_
timestamp 1635444444
transform 1 0 2392 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_79_30
timestamp 1635444444
transform 1 0 3864 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1635444444
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1635444444
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_42
timestamp 1635444444
transform 1 0 4968 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1635444444
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_54
timestamp 1635444444
transform 1 0 6072 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1635444444
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1635444444
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1635444444
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1635444444
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1635444444
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1635444444
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1635444444
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1635444444
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1635444444
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1635444444
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_93
timestamp 1635444444
transform 1 0 9660 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_99
timestamp 1635444444
transform 1 0 10212 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_97
timestamp 1635444444
transform 1 0 10028 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635444444
transform 1 0 9936 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1635444444
transform -1 0 10856 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1635444444
transform -1 0 10856 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_7
timestamp 1635444444
transform 1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1635444444
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1635444444
transform -1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1635444444
transform -1 0 2484 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_15
timestamp 1635444444
transform 1 0 2484 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_23
timestamp 1635444444
transform 1 0 3220 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1635444444
transform 1 0 2852 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_30
timestamp 1635444444
transform 1 0 3864 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _182_
timestamp 1635444444
transform 1 0 3588 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_42
timestamp 1635444444
transform 1 0 4968 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1635444444
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1635444444
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1635444444
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1635444444
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1635444444
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_93
timestamp 1635444444
transform 1 0 9660 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_99
timestamp 1635444444
transform 1 0 10212 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635444444
transform 1 0 9936 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1635444444
transform -1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_7
timestamp 1635444444
transform 1 0 1748 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1635444444
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1635444444
transform -1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_18
timestamp 1635444444
transform 1 0 2760 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _181_
timestamp 1635444444
transform 1 0 2484 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_26
timestamp 1635444444
transform 1 0 3496 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_32
timestamp 1635444444
transform 1 0 4048 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1635444444
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _184_
timestamp 1635444444
transform 1 0 3772 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_44
timestamp 1635444444
transform 1 0 5152 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_56
timestamp 1635444444
transform 1 0 6256 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_68
timestamp 1635444444
transform 1 0 7360 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_80
timestamp 1635444444
transform 1 0 8464 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1635444444
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1635444444
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_97
timestamp 1635444444
transform 1 0 10028 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1635444444
transform -1 0 10856 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_7
timestamp 1635444444
transform 1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1635444444
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1635444444
transform -1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1635444444
transform -1 0 2484 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_15
timestamp 1635444444
transform 1 0 2484 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_22
timestamp 1635444444
transform 1 0 3128 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _183_
timestamp 1635444444
transform 1 0 2852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_34
timestamp 1635444444
transform 1 0 4232 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_46
timestamp 1635444444
transform 1 0 5336 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_54
timestamp 1635444444
transform 1 0 6072 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1635444444
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1635444444
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1635444444
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1635444444
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_93
timestamp 1635444444
transform 1 0 9660 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_99
timestamp 1635444444
transform 1 0 10212 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1635444444
transform 1 0 9936 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1635444444
transform -1 0 10856 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_84_7
timestamp 1635444444
transform 1 0 1748 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1635444444
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1635444444
transform -1 0 1748 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_18
timestamp 1635444444
transform 1 0 2760 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _185_
timestamp 1635444444
transform 1 0 2484 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_84_26
timestamp 1635444444
transform 1 0 3496 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1635444444
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1635444444
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1635444444
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1635444444
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1635444444
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1635444444
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1635444444
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_85
timestamp 1635444444
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1635444444
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_97
timestamp 1635444444
transform 1 0 10028 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1635444444
transform -1 0 10856 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_7
timestamp 1635444444
transform 1 0 1748 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_7
timestamp 1635444444
transform 1 0 1748 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1635444444
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1635444444
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1635444444
transform -1 0 1748 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1635444444
transform -1 0 1748 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1635444444
transform -1 0 2484 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1635444444
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_13
timestamp 1635444444
transform 1 0 2300 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_17
timestamp 1635444444
transform 1 0 2668 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_24
timestamp 1635444444
transform 1 0 3312 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _187_
timestamp 1635444444
transform -1 0 2668 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _190_
timestamp 1635444444
transform 1 0 3036 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1635444444
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1635444444
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _180_
timestamp 1635444444
transform 1 0 3772 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1635444444
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1635444444
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_39
timestamp 1635444444
transform 1 0 4692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_51
timestamp 1635444444
transform 1 0 5796 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1635444444
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1635444444
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_63
timestamp 1635444444
transform 1 0 6900 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1635444444
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1635444444
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_75
timestamp 1635444444
transform 1 0 8004 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1635444444
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1635444444
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_85
timestamp 1635444444
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1635444444
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_93
timestamp 1635444444
transform 1 0 9660 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_99
timestamp 1635444444
transform 1 0 10212 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_97
timestamp 1635444444
transform 1 0 10028 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1635444444
transform 1 0 9936 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1635444444
transform -1 0 10856 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1635444444
transform -1 0 10856 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_7
timestamp 1635444444
transform 1 0 1748 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1635444444
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1635444444
transform -1 0 1748 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1635444444
transform -1 0 2484 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_15
timestamp 1635444444
transform 1 0 2484 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_22
timestamp 1635444444
transform 1 0 3128 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _188_
timestamp 1635444444
transform -1 0 3128 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_29
timestamp 1635444444
transform 1 0 3772 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _189_
timestamp 1635444444
transform 1 0 3496 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_41
timestamp 1635444444
transform 1 0 4876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_53
timestamp 1635444444
transform 1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1635444444
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1635444444
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1635444444
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1635444444
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_93
timestamp 1635444444
transform 1 0 9660 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_99
timestamp 1635444444
transform 1 0 10212 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1635444444
transform 1 0 9936 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1635444444
transform -1 0 10856 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_10
timestamp 1635444444
transform 1 0 2024 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1635444444
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _239_
timestamp 1635444444
transform -1 0 2024 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_88_18
timestamp 1635444444
transform 1 0 2760 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1635444444
transform -1 0 2760 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1635444444
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1635444444
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _186_
timestamp 1635444444
transform 1 0 3772 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_88_39
timestamp 1635444444
transform 1 0 4692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_51
timestamp 1635444444
transform 1 0 5796 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_63
timestamp 1635444444
transform 1 0 6900 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_75
timestamp 1635444444
transform 1 0 8004 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1635444444
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_85
timestamp 1635444444
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1635444444
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_97
timestamp 1635444444
transform 1 0 10028 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1635444444
transform -1 0 10856 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_89_3
timestamp 1635444444
transform 1 0 1380 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1635444444
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _238_
timestamp 1635444444
transform 1 0 1932 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_89_19
timestamp 1635444444
transform 1 0 2852 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1635444444
transform 1 0 3220 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_27
timestamp 1635444444
transform 1 0 3588 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_34
timestamp 1635444444
transform 1 0 4232 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _191_
timestamp 1635444444
transform 1 0 3956 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_89_46
timestamp 1635444444
transform 1 0 5336 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_54
timestamp 1635444444
transform 1 0 6072 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1635444444
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1635444444
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1635444444
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1635444444
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_93
timestamp 1635444444
transform 1 0 9660 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_99
timestamp 1635444444
transform 1 0 10212 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1635444444
transform 1 0 9936 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1635444444
transform -1 0 10856 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_90_10
timestamp 1635444444
transform 1 0 2024 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1635444444
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _240_
timestamp 1635444444
transform 1 0 1380 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_90_21
timestamp 1635444444
transform 1 0 3036 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _241_
timestamp 1635444444
transform -1 0 3036 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1635444444
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_33
timestamp 1635444444
transform 1 0 4140 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1635444444
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1635444444
transform 1 0 3772 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_45
timestamp 1635444444
transform 1 0 5244 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_57
timestamp 1635444444
transform 1 0 6348 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_69
timestamp 1635444444
transform 1 0 7452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1635444444
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_85
timestamp 1635444444
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1635444444
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_97
timestamp 1635444444
transform 1 0 10028 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1635444444
transform -1 0 10856 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_91_3
timestamp 1635444444
transform 1 0 1380 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1635444444
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _237_
timestamp 1635444444
transform -1 0 2576 0 -1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_91_16
timestamp 1635444444
transform 1 0 2576 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _179_
timestamp 1635444444
transform 1 0 2944 0 -1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_91_30
timestamp 1635444444
transform 1 0 3864 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_42
timestamp 1635444444
transform 1 0 4968 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_54
timestamp 1635444444
transform 1 0 6072 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1635444444
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1635444444
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1635444444
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1635444444
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_93
timestamp 1635444444
transform 1 0 9660 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_99
timestamp 1635444444
transform 1 0 10212 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1635444444
transform 1 0 9936 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1635444444
transform -1 0 10856 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_92_10
timestamp 1635444444
transform 1 0 2024 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_10
timestamp 1635444444
transform 1 0 2024 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1635444444
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1635444444
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _242_
timestamp 1635444444
transform -1 0 2024 0 1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _243_
timestamp 1635444444
transform 1 0 1380 0 -1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_92_20
timestamp 1635444444
transform 1 0 2944 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_18
timestamp 1635444444
transform 1 0 2760 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_25
timestamp 1635444444
transform 1 0 3404 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _223_
timestamp 1635444444
transform -1 0 3404 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _230_
timestamp 1635444444
transform 1 0 2576 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1635444444
transform -1 0 2760 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_32
timestamp 1635444444
transform 1 0 4048 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_37
timestamp 1635444444
transform 1 0 4508 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1635444444
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _224_
timestamp 1635444444
transform 1 0 3772 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_44
timestamp 1635444444
transform 1 0 5152 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_49
timestamp 1635444444
transform 1 0 5612 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_92_56
timestamp 1635444444
transform 1 0 6256 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1635444444
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1635444444
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1635444444
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_68
timestamp 1635444444
transform 1 0 7360 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1635444444
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_80
timestamp 1635444444
transform 1 0 8464 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_85
timestamp 1635444444
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_81
timestamp 1635444444
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1635444444
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_97
timestamp 1635444444
transform 1 0 10028 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_93_93
timestamp 1635444444
transform 1 0 9660 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_99
timestamp 1635444444
transform 1 0 10212 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1635444444
transform 1 0 9936 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1635444444
transform -1 0 10856 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1635444444
transform -1 0 10856 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_7
timestamp 1635444444
transform 1 0 1748 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1635444444
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1635444444
transform -1 0 1748 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1635444444
transform 1 0 2116 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_15
timestamp 1635444444
transform 1 0 2484 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_22
timestamp 1635444444
transform 1 0 3128 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _225_
timestamp 1635444444
transform 1 0 2852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1635444444
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1635444444
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1635444444
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1635444444
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1635444444
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1635444444
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1635444444
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_85
timestamp 1635444444
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1635444444
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_97
timestamp 1635444444
transform 1 0 10028 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1635444444
transform -1 0 10856 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_7
timestamp 1635444444
transform 1 0 1748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1635444444
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1635444444
transform -1 0 1748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1635444444
transform -1 0 2484 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1635444444
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1635444444
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_39
timestamp 1635444444
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1635444444
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1635444444
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1635444444
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1635444444
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1635444444
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1635444444
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_93
timestamp 1635444444
transform 1 0 9660 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_99
timestamp 1635444444
transform 1 0 10212 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1635444444
transform 1 0 9936 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1635444444
transform -1 0 10856 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_7
timestamp 1635444444
transform 1 0 1748 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1635444444
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1635444444
transform -1 0 1748 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_19
timestamp 1635444444
transform 1 0 2852 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1635444444
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1635444444
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1635444444
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1635444444
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1635444444
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1635444444
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1635444444
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1635444444
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_85
timestamp 1635444444
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1635444444
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_97
timestamp 1635444444
transform 1 0 10028 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1635444444
transform -1 0 10856 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_7
timestamp 1635444444
transform 1 0 1748 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1635444444
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1635444444
transform -1 0 1748 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1635444444
transform -1 0 2484 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1635444444
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1635444444
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1635444444
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1635444444
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1635444444
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1635444444
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1635444444
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1635444444
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1635444444
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_93
timestamp 1635444444
transform 1 0 9660 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_99
timestamp 1635444444
transform 1 0 10212 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1635444444
transform 1 0 9936 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1635444444
transform -1 0 10856 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_7
timestamp 1635444444
transform 1 0 1748 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1635444444
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1635444444
transform -1 0 1748 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_19
timestamp 1635444444
transform 1 0 2852 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1635444444
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_29
timestamp 1635444444
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1635444444
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_41
timestamp 1635444444
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_53
timestamp 1635444444
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_65
timestamp 1635444444
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1635444444
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1635444444
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_85
timestamp 1635444444
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1635444444
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_97
timestamp 1635444444
transform 1 0 10028 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1635444444
transform -1 0 10856 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_10
timestamp 1635444444
transform 1 0 2024 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_7
timestamp 1635444444
transform 1 0 1748 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1635444444
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1635444444
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _247_
timestamp 1635444444
transform -1 0 2024 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1635444444
transform -1 0 1748 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1635444444
transform 1 0 2116 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_18
timestamp 1635444444
transform 1 0 2760 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_15
timestamp 1635444444
transform 1 0 2484 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_19
timestamp 1635444444
transform 1 0 2852 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_23
timestamp 1635444444
transform 1 0 3220 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1635444444
transform 1 0 2944 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1635444444
transform -1 0 2760 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_26
timestamp 1635444444
transform 1 0 3496 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_29
timestamp 1635444444
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_35
timestamp 1635444444
transform 1 0 4324 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1635444444
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_41
timestamp 1635444444
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_47
timestamp 1635444444
transform 1 0 5428 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_53
timestamp 1635444444
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1635444444
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1635444444
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1635444444
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_65
timestamp 1635444444
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1635444444
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1635444444
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1635444444
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_85
timestamp 1635444444
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1635444444
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1635444444
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_97
timestamp 1635444444
transform 1 0 10028 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_99_93
timestamp 1635444444
transform 1 0 9660 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_99
timestamp 1635444444
transform 1 0 10212 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635444444
transform 1 0 9936 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1635444444
transform -1 0 10856 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1635444444
transform -1 0 10856 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_10
timestamp 1635444444
transform 1 0 2024 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1635444444
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _246_
timestamp 1635444444
transform 1 0 1380 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_101_24
timestamp 1635444444
transform 1 0 3312 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _245_
timestamp 1635444444
transform 1 0 2392 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_101_32
timestamp 1635444444
transform 1 0 4048 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1635444444
transform 1 0 3680 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_44
timestamp 1635444444
transform 1 0 5152 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1635444444
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1635444444
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1635444444
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_81
timestamp 1635444444
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_93
timestamp 1635444444
transform 1 0 9660 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_99
timestamp 1635444444
transform 1 0 10212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635444444
transform 1 0 9936 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1635444444
transform -1 0 10856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_102_10
timestamp 1635444444
transform 1 0 2024 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1635444444
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _248_
timestamp 1635444444
transform 1 0 1380 0 1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_102_24
timestamp 1635444444
transform 1 0 3312 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _244_
timestamp 1635444444
transform 1 0 2392 0 1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_102_29
timestamp 1635444444
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1635444444
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_41
timestamp 1635444444
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_53
timestamp 1635444444
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1635444444
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1635444444
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1635444444
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_85
timestamp 1635444444
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1635444444
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_97
timestamp 1635444444
transform 1 0 10028 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1635444444
transform -1 0 10856 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_103_10
timestamp 1635444444
transform 1 0 2024 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1635444444
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _249_
timestamp 1635444444
transform -1 0 2024 0 -1 58752
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_103_18
timestamp 1635444444
transform 1 0 2760 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1635444444
transform -1 0 2760 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_30
timestamp 1635444444
transform 1 0 3864 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_42
timestamp 1635444444
transform 1 0 4968 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_54
timestamp 1635444444
transform 1 0 6072 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1635444444
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1635444444
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1635444444
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_81
timestamp 1635444444
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_93
timestamp 1635444444
transform 1 0 9660 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_103_99
timestamp 1635444444
transform 1 0 10212 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1635444444
transform 1 0 9936 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1635444444
transform -1 0 10856 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_10
timestamp 1635444444
transform 1 0 2024 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1635444444
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _250_
timestamp 1635444444
transform -1 0 2024 0 1 58752
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_104_18
timestamp 1635444444
transform 1 0 2760 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1635444444
transform -1 0 2760 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_104_26
timestamp 1635444444
transform 1 0 3496 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1635444444
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1635444444
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_41
timestamp 1635444444
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_53
timestamp 1635444444
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_65
timestamp 1635444444
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1635444444
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1635444444
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_85
timestamp 1635444444
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1635444444
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_104_97
timestamp 1635444444
transform 1 0 10028 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1635444444
transform -1 0 10856 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_7
timestamp 1635444444
transform 1 0 1748 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_7
timestamp 1635444444
transform 1 0 1748 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1635444444
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1635444444
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1635444444
transform -1 0 1748 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1635444444
transform -1 0 1748 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1635444444
transform -1 0 2484 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1635444444
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_19
timestamp 1635444444
transform 1 0 2852 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1635444444
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1635444444
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1635444444
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1635444444
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_39
timestamp 1635444444
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1635444444
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1635444444
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1635444444
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1635444444
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1635444444
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1635444444
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1635444444
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_65
timestamp 1635444444
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1635444444
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_105_81
timestamp 1635444444
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1635444444
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_85
timestamp 1635444444
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1635444444
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_105_93
timestamp 1635444444
transform 1 0 9660 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_99
timestamp 1635444444
transform 1 0 10212 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_97
timestamp 1635444444
transform 1 0 10028 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1635444444
transform 1 0 9936 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1635444444
transform -1 0 10856 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1635444444
transform -1 0 10856 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_7
timestamp 1635444444
transform 1 0 1748 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1635444444
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1635444444
transform -1 0 1748 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_19
timestamp 1635444444
transform 1 0 2852 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_31
timestamp 1635444444
transform 1 0 3956 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_43
timestamp 1635444444
transform 1 0 5060 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1635444444
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1635444444
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1635444444
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1635444444
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_81
timestamp 1635444444
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_93
timestamp 1635444444
transform 1 0 9660 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_99
timestamp 1635444444
transform 1 0 10212 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635444444
transform 1 0 9936 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1635444444
transform -1 0 10856 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_7
timestamp 1635444444
transform 1 0 1748 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1635444444
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1635444444
transform -1 0 1748 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1635444444
transform -1 0 2484 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_108_15
timestamp 1635444444
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1635444444
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_29
timestamp 1635444444
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1635444444
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_41
timestamp 1635444444
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_53
timestamp 1635444444
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_65
timestamp 1635444444
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1635444444
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1635444444
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_85
timestamp 1635444444
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1635444444
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_97
timestamp 1635444444
transform 1 0 10028 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1635444444
transform -1 0 10856 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_109_7
timestamp 1635444444
transform 1 0 1748 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1635444444
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _254_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2852 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1635444444
transform -1 0 1748 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_109_19
timestamp 1635444444
transform 1 0 2852 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_31
timestamp 1635444444
transform 1 0 3956 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_43
timestamp 1635444444
transform 1 0 5060 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1635444444
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1635444444
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1635444444
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1635444444
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_81
timestamp 1635444444
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_109_93
timestamp 1635444444
transform 1 0 9660 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_109_99
timestamp 1635444444
transform 1 0 10212 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1635444444
transform 1 0 9936 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1635444444
transform -1 0 10856 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_110_7
timestamp 1635444444
transform 1 0 1748 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1635444444
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _253_
timestamp 1635444444
transform -1 0 2852 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1635444444
transform -1 0 1748 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_110_19
timestamp 1635444444
transform 1 0 2852 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1635444444
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1635444444
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1635444444
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1635444444
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1635444444
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_65
timestamp 1635444444
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1635444444
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1635444444
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_85
timestamp 1635444444
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1635444444
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_110_97
timestamp 1635444444
transform 1 0 10028 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1635444444
transform -1 0 10856 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_111_3
timestamp 1635444444
transform 1 0 1380 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1635444444
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _255_
timestamp 1635444444
transform -1 0 2300 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_111_13
timestamp 1635444444
transform 1 0 2300 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _252_
timestamp 1635444444
transform 1 0 2668 0 -1 63104
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_111_27
timestamp 1635444444
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_39
timestamp 1635444444
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1635444444
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1635444444
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_57
timestamp 1635444444
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1635444444
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_69
timestamp 1635444444
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_81
timestamp 1635444444
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_93
timestamp 1635444444
transform 1 0 9660 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_111_99
timestamp 1635444444
transform 1 0 10212 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1635444444
transform 1 0 9936 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1635444444
transform -1 0 10856 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_112_7
timestamp 1635444444
transform 1 0 1748 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_113_7
timestamp 1635444444
transform 1 0 1748 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1635444444
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1635444444
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _256_
timestamp 1635444444
transform -1 0 2852 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1635444444
transform -1 0 1748 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1635444444
transform -1 0 1748 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_112_13
timestamp 1635444444
transform 1 0 2300 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_112_24
timestamp 1635444444
transform 1 0 3312 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_113_19
timestamp 1635444444
transform 1 0 2852 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _251_
timestamp 1635444444
transform 1 0 2392 0 1 63104
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_112_33
timestamp 1635444444
transform 1 0 4140 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_31
timestamp 1635444444
transform 1 0 3956 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1635444444
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1635444444
transform 1 0 3772 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_112_45
timestamp 1635444444
transform 1 0 5244 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_43
timestamp 1635444444
transform 1 0 5060 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_57
timestamp 1635444444
transform 1 0 6348 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1635444444
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1635444444
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1635444444
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_69
timestamp 1635444444
transform 1 0 7452 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1635444444
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_112_81
timestamp 1635444444
transform 1 0 8556 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_85
timestamp 1635444444
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_81
timestamp 1635444444
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1635444444
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_112_97
timestamp 1635444444
transform 1 0 10028 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_113_93
timestamp 1635444444
transform 1 0 9660 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_113_99
timestamp 1635444444
transform 1 0 10212 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1635444444
transform 1 0 9936 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1635444444
transform -1 0 10856 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1635444444
transform -1 0 10856 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_114_3
timestamp 1635444444
transform 1 0 1380 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_9
timestamp 1635444444
transform 1 0 1932 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1635444444
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _257_
timestamp 1635444444
transform -1 0 2760 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_114_18
timestamp 1635444444
transform 1 0 2760 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_114_26
timestamp 1635444444
transform 1 0 3496 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_114_33
timestamp 1635444444
transform 1 0 4140 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1635444444
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1635444444
transform 1 0 3772 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_114_45
timestamp 1635444444
transform 1 0 5244 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_57
timestamp 1635444444
transform 1 0 6348 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_69
timestamp 1635444444
transform 1 0 7452 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_114_81
timestamp 1635444444
transform 1 0 8556 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_114_85
timestamp 1635444444
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1635444444
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_114_97
timestamp 1635444444
transform 1 0 10028 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1635444444
transform -1 0 10856 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_115_7
timestamp 1635444444
transform 1 0 1748 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1635444444
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1635444444
transform -1 0 1748 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_115_15
timestamp 1635444444
transform 1 0 2484 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_22
timestamp 1635444444
transform 1 0 3128 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _227_
timestamp 1635444444
transform 1 0 2760 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_115_34
timestamp 1635444444
transform 1 0 4232 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_46
timestamp 1635444444
transform 1 0 5336 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_115_54
timestamp 1635444444
transform 1 0 6072 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_115_57
timestamp 1635444444
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1635444444
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_69
timestamp 1635444444
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_81
timestamp 1635444444
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_115_93
timestamp 1635444444
transform 1 0 9660 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_99
timestamp 1635444444
transform 1 0 10212 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1635444444
transform 1 0 9936 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1635444444
transform -1 0 10856 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_116_11
timestamp 1635444444
transform 1 0 2116 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_3
timestamp 1635444444
transform 1 0 1380 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1635444444
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1635444444
transform -1 0 2116 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_116_19
timestamp 1635444444
transform 1 0 2852 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1635444444
transform -1 0 2852 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1635444444
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_29
timestamp 1635444444
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1635444444
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_41
timestamp 1635444444
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_53
timestamp 1635444444
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_65
timestamp 1635444444
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_77
timestamp 1635444444
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1635444444
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_85
timestamp 1635444444
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1635444444
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_116_97
timestamp 1635444444
transform 1 0 10028 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1635444444
transform -1 0 10856 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_117_11
timestamp 1635444444
transform 1 0 2116 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_117_3
timestamp 1635444444
transform 1 0 1380 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1635444444
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1635444444
transform -1 0 2116 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_117_23
timestamp 1635444444
transform 1 0 3220 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1635444444
transform 1 0 2852 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_117_35
timestamp 1635444444
transform 1 0 4324 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_47
timestamp 1635444444
transform 1 0 5428 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_55
timestamp 1635444444
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1635444444
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1635444444
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1635444444
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_81
timestamp 1635444444
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_93
timestamp 1635444444
transform 1 0 9660 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_99
timestamp 1635444444
transform 1 0 10212 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635444444
transform 1 0 9936 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1635444444
transform -1 0 10856 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_118_11
timestamp 1635444444
transform 1 0 2116 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_3
timestamp 1635444444
transform 1 0 1380 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1635444444
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1635444444
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1635444444
transform -1 0 2116 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1635444444
transform 1 0 1380 0 -1 67456
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_118_19
timestamp 1635444444
transform 1 0 2852 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_13
timestamp 1635444444
transform 1 0 2300 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_25
timestamp 1635444444
transform 1 0 3404 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1635444444
transform -1 0 2852 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1635444444
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_29
timestamp 1635444444
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_37
timestamp 1635444444
transform 1 0 4508 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1635444444
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_41
timestamp 1635444444
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_49
timestamp 1635444444
transform 1 0 5612 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_118_53
timestamp 1635444444
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1635444444
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1635444444
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1635444444
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_65
timestamp 1635444444
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1635444444
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_119_69
timestamp 1635444444
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1635444444
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_85
timestamp 1635444444
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_81
timestamp 1635444444
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1635444444
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_118_97
timestamp 1635444444
transform 1 0 10028 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_119_101
timestamp 1635444444
transform 1 0 10396 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_119_93
timestamp 1635444444
transform 1 0 9660 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1635444444
transform -1 0 10856 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1635444444
transform -1 0 10856 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_120_3
timestamp 1635444444
transform 1 0 1380 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_120_9
timestamp 1635444444
transform 1 0 1932 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1635444444
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1635444444
transform 1 0 1564 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_120_23
timestamp 1635444444
transform 1 0 3220 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _259_
timestamp 1635444444
transform -1 0 3220 0 1 67456
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1635444444
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_29
timestamp 1635444444
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1635444444
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_41
timestamp 1635444444
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_53
timestamp 1635444444
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_65
timestamp 1635444444
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1635444444
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1635444444
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_85
timestamp 1635444444
transform 1 0 8924 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1635444444
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_120_93
timestamp 1635444444
transform 1 0 9660 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_99
timestamp 1635444444
transform 1 0 10212 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635444444
transform 1 0 9936 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1635444444
transform -1 0 10856 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_11
timestamp 1635444444
transform 1 0 2116 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1635444444
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _260_
timestamp 1635444444
transform -1 0 2116 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_121_15
timestamp 1635444444
transform 1 0 2484 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _258_
timestamp 1635444444
transform 1 0 2576 0 -1 68544
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_121_26
timestamp 1635444444
transform 1 0 3496 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_38
timestamp 1635444444
transform 1 0 4600 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _261_
timestamp 1635444444
transform -1 0 4600 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_121_50
timestamp 1635444444
transform 1 0 5704 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1635444444
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1635444444
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1635444444
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_81
timestamp 1635444444
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_101
timestamp 1635444444
transform 1 0 10396 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_121_93
timestamp 1635444444
transform 1 0 9660 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1635444444
transform -1 0 10856 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1635444444
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1635444444
transform 1 0 1380 0 1 68544
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_122_13
timestamp 1635444444
transform 1 0 2300 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_122_25
timestamp 1635444444
transform 1 0 3404 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_122_37
timestamp 1635444444
transform 1 0 4508 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1635444444
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_2  _262_
timestamp 1635444444
transform -1 0 4508 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_49
timestamp 1635444444
transform 1 0 5612 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_61
timestamp 1635444444
transform 1 0 6716 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_73
timestamp 1635444444
transform 1 0 7820 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_81
timestamp 1635444444
transform 1 0 8556 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_122_85
timestamp 1635444444
transform 1 0 8924 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1635444444
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_122_93
timestamp 1635444444
transform 1 0 9660 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_99
timestamp 1635444444
transform 1 0 10212 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635444444
transform 1 0 9936 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1635444444
transform -1 0 10856 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1635444444
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1635444444
transform 1 0 1380 0 -1 69632
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_123_13
timestamp 1635444444
transform 1 0 2300 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _265_
timestamp 1635444444
transform 1 0 2852 0 -1 69632
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_123_29
timestamp 1635444444
transform 1 0 3772 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _266_
timestamp 1635444444
transform 1 0 4140 0 -1 69632
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_123_43
timestamp 1635444444
transform 1 0 5060 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1635444444
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_57
timestamp 1635444444
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1635444444
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_69
timestamp 1635444444
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_81
timestamp 1635444444
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_101
timestamp 1635444444
transform 1 0 10396 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_123_93
timestamp 1635444444
transform 1 0 9660 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1635444444
transform -1 0 10856 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1635444444
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1635444444
transform 1 0 1380 0 1 69632
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_124_13
timestamp 1635444444
transform 1 0 2300 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_124_20
timestamp 1635444444
transform 1 0 2944 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1635444444
transform 1 0 2668 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_124_29
timestamp 1635444444
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1635444444
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_41
timestamp 1635444444
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_53
timestamp 1635444444
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_65
timestamp 1635444444
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1635444444
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1635444444
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_85
timestamp 1635444444
transform 1 0 8924 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1635444444
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_124_93
timestamp 1635444444
transform 1 0 9660 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_124_99
timestamp 1635444444
transform 1 0 10212 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635444444
transform 1 0 9936 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1635444444
transform -1 0 10856 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_126_11
timestamp 1635444444
transform 1 0 2116 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1635444444
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1635444444
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _263_
timestamp 1635444444
transform 1 0 1380 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1635444444
transform 1 0 1380 0 -1 70720
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_125_13
timestamp 1635444444
transform 1 0 2300 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_125_25
timestamp 1635444444
transform 1 0 3404 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_18
timestamp 1635444444
transform 1 0 2760 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _264_
timestamp 1635444444
transform 1 0 2668 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1635444444
transform 1 0 2484 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_37
timestamp 1635444444
transform 1 0 4508 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_126_26
timestamp 1635444444
transform 1 0 3496 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_126_29
timestamp 1635444444
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1635444444
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_125_49
timestamp 1635444444
transform 1 0 5612 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_126_41
timestamp 1635444444
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1635444444
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_57
timestamp 1635444444
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_53
timestamp 1635444444
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1635444444
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_69
timestamp 1635444444
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_65
timestamp 1635444444
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1635444444
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_125_81
timestamp 1635444444
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1635444444
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_126_85
timestamp 1635444444
transform 1 0 8924 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1635444444
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_125_101
timestamp 1635444444
transform 1 0 10396 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_125_93
timestamp 1635444444
transform 1 0 9660 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_126_93
timestamp 1635444444
transform 1 0 9660 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_126_99
timestamp 1635444444
transform 1 0 10212 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1635444444
transform 1 0 9936 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1635444444
transform -1 0 10856 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1635444444
transform -1 0 10856 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_127_10
timestamp 1635444444
transform 1 0 2024 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_127_6
timestamp 1635444444
transform 1 0 1656 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1635444444
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _267_
timestamp 1635444444
transform -1 0 2852 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1635444444
transform -1 0 1656 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_127_19
timestamp 1635444444
transform 1 0 2852 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_31
timestamp 1635444444
transform 1 0 3956 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_43
timestamp 1635444444
transform 1 0 5060 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1635444444
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_57
timestamp 1635444444
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1635444444
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_69
timestamp 1635444444
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_81
timestamp 1635444444
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_101
timestamp 1635444444
transform 1 0 10396 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_127_93
timestamp 1635444444
transform 1 0 9660 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1635444444
transform -1 0 10856 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_128_10
timestamp 1635444444
transform 1 0 2024 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_128_6
timestamp 1635444444
transform 1 0 1656 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1635444444
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _268_
timestamp 1635444444
transform -1 0 2852 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1635444444
transform -1 0 1656 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_128_19
timestamp 1635444444
transform 1 0 2852 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 1635444444
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_29
timestamp 1635444444
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1635444444
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_41
timestamp 1635444444
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_53
timestamp 1635444444
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_65
timestamp 1635444444
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1635444444
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1635444444
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_85
timestamp 1635444444
transform 1 0 8924 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1635444444
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_128_93
timestamp 1635444444
transform 1 0 9660 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_128_99
timestamp 1635444444
transform 1 0 10212 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1635444444
transform 1 0 9936 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1635444444
transform -1 0 10856 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_129_6
timestamp 1635444444
transform 1 0 1656 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1635444444
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1635444444
transform -1 0 1656 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1635444444
transform -1 0 2300 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_129_13
timestamp 1635444444
transform 1 0 2300 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_25
timestamp 1635444444
transform 1 0 3404 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_37
timestamp 1635444444
transform 1 0 4508 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_49
timestamp 1635444444
transform 1 0 5612 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1635444444
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_57
timestamp 1635444444
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1635444444
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_69
timestamp 1635444444
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_81
timestamp 1635444444
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_101
timestamp 1635444444
transform 1 0 10396 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_129_93
timestamp 1635444444
transform 1 0 9660 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1635444444
transform -1 0 10856 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_130_10
timestamp 1635444444
transform 1 0 2024 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_130_6
timestamp 1635444444
transform 1 0 1656 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1635444444
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _269_
timestamp 1635444444
transform -1 0 2852 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1635444444
transform -1 0 1656 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_130_19
timestamp 1635444444
transform 1 0 2852 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 1635444444
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_29
timestamp 1635444444
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1635444444
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_41
timestamp 1635444444
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_53
timestamp 1635444444
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_65
timestamp 1635444444
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1635444444
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1635444444
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_85
timestamp 1635444444
transform 1 0 8924 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1635444444
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_130_93
timestamp 1635444444
transform 1 0 9660 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_130_99
timestamp 1635444444
transform 1 0 10212 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1635444444
transform 1 0 9936 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1635444444
transform -1 0 10856 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_131_10
timestamp 1635444444
transform 1 0 2024 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_131_6
timestamp 1635444444
transform 1 0 1656 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1635444444
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _270_
timestamp 1635444444
transform -1 0 2852 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1635444444
transform -1 0 1656 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_19
timestamp 1635444444
transform 1 0 2852 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_31
timestamp 1635444444
transform 1 0 3956 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_43
timestamp 1635444444
transform 1 0 5060 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_131_55
timestamp 1635444444
transform 1 0 6164 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_57
timestamp 1635444444
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1635444444
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_69
timestamp 1635444444
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_81
timestamp 1635444444
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_101
timestamp 1635444444
transform 1 0 10396 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_131_93
timestamp 1635444444
transform 1 0 9660 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1635444444
transform -1 0 10856 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_132_10
timestamp 1635444444
transform 1 0 2024 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_132_6
timestamp 1635444444
transform 1 0 1656 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_133_3
timestamp 1635444444
transform 1 0 1380 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1635444444
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1635444444
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _271_
timestamp 1635444444
transform -1 0 2852 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _272_
timestamp 1635444444
transform -1 0 2392 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1635444444
transform -1 0 1656 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_132_19
timestamp 1635444444
transform 1 0 2852 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_133_14
timestamp 1635444444
transform 1 0 2392 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _274_
timestamp 1635444444
transform -1 0 3496 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1635444444
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_32
timestamp 1635444444
transform 1 0 4048 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_26
timestamp 1635444444
transform 1 0 3496 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_38
timestamp 1635444444
transform 1 0 4600 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1635444444
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1635444444
transform 1 0 3772 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_44
timestamp 1635444444
transform 1 0 5152 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_50
timestamp 1635444444
transform 1 0 5704 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_132_56
timestamp 1635444444
transform 1 0 6256 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_57
timestamp 1635444444
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1635444444
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_68
timestamp 1635444444
transform 1 0 7360 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_69
timestamp 1635444444
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_132_80
timestamp 1635444444
transform 1 0 8464 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_132_85
timestamp 1635444444
transform 1 0 8924 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_81
timestamp 1635444444
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1635444444
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_132_93
timestamp 1635444444
transform 1 0 9660 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_99
timestamp 1635444444
transform 1 0 10212 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_133_101
timestamp 1635444444
transform 1 0 10396 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_133_93
timestamp 1635444444
transform 1 0 9660 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1635444444
transform 1 0 9936 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1635444444
transform -1 0 10856 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1635444444
transform -1 0 10856 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_134_3
timestamp 1635444444
transform 1 0 1380 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1635444444
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _273_
timestamp 1635444444
transform -1 0 2392 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_134_14
timestamp 1635444444
transform 1 0 2392 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_134_21
timestamp 1635444444
transform 1 0 3036 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1635444444
transform -1 0 3036 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1635444444
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_29
timestamp 1635444444
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1635444444
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_41
timestamp 1635444444
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_53
timestamp 1635444444
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_65
timestamp 1635444444
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1635444444
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1635444444
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_85
timestamp 1635444444
transform 1 0 8924 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1635444444
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_134_93
timestamp 1635444444
transform 1 0 9660 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_99
timestamp 1635444444
transform 1 0 10212 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1635444444
transform 1 0 9936 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1635444444
transform -1 0 10856 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_135_6
timestamp 1635444444
transform 1 0 1656 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1635444444
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1635444444
transform -1 0 1656 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1635444444
transform 1 0 2024 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_13
timestamp 1635444444
transform 1 0 2300 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_25
timestamp 1635444444
transform 1 0 3404 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_37
timestamp 1635444444
transform 1 0 4508 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_49
timestamp 1635444444
transform 1 0 5612 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_55
timestamp 1635444444
transform 1 0 6164 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_57
timestamp 1635444444
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1635444444
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_69
timestamp 1635444444
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_81
timestamp 1635444444
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_135_101
timestamp 1635444444
transform 1 0 10396 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_135_93
timestamp 1635444444
transform 1 0 9660 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1635444444
transform -1 0 10856 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_6
timestamp 1635444444
transform 1 0 1656 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1635444444
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1635444444
transform -1 0 1656 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1635444444
transform 1 0 2024 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_13
timestamp 1635444444
transform 1 0 2300 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_136_20
timestamp 1635444444
transform 1 0 2944 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1635444444
transform -1 0 2944 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_136_29
timestamp 1635444444
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1635444444
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_41
timestamp 1635444444
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_53
timestamp 1635444444
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_65
timestamp 1635444444
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1635444444
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1635444444
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_85
timestamp 1635444444
transform 1 0 8924 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1635444444
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_136_93
timestamp 1635444444
transform 1 0 9660 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_99
timestamp 1635444444
transform 1 0 10212 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1635444444
transform 1 0 9936 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1635444444
transform -1 0 10856 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_6
timestamp 1635444444
transform 1 0 1656 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1635444444
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1635444444
transform -1 0 1656 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1635444444
transform -1 0 2300 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_13
timestamp 1635444444
transform 1 0 2300 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_137_20
timestamp 1635444444
transform 1 0 2944 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1635444444
transform 1 0 2668 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_137_32
timestamp 1635444444
transform 1 0 4048 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_44
timestamp 1635444444
transform 1 0 5152 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_57
timestamp 1635444444
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1635444444
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_69
timestamp 1635444444
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_81
timestamp 1635444444
transform 1 0 8556 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_137_93
timestamp 1635444444
transform 1 0 9660 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_99
timestamp 1635444444
transform 1 0 10212 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1635444444
transform 1 0 9936 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1635444444
transform -1 0 10856 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_6
timestamp 1635444444
transform 1 0 1656 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1635444444
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1635444444
transform -1 0 1656 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1635444444
transform -1 0 2300 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_13
timestamp 1635444444
transform 1 0 2300 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_138_20
timestamp 1635444444
transform 1 0 2944 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1635444444
transform 1 0 2668 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_32
timestamp 1635444444
transform 1 0 4048 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1635444444
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1635444444
transform 1 0 3772 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_44
timestamp 1635444444
transform 1 0 5152 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_57
timestamp 1635444444
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1635444444
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_69
timestamp 1635444444
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1635444444
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_85
timestamp 1635444444
transform 1 0 8924 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1635444444
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1635444444
transform 1 0 9292 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_92
timestamp 1635444444
transform 1 0 9568 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_99
timestamp 1635444444
transform 1 0 10212 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1635444444
transform 1 0 9936 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1635444444
transform -1 0 10856 0 1 77248
box -38 -48 314 592
<< labels >>
rlabel metal4 s 2575 2128 2895 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 5839 2128 6159 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 9103 2128 9423 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 4207 2128 4527 77840 6 vssd1
port 1 nsew ground input
rlabel metal4 s 7471 2128 7791 77840 6 vssd1
port 1 nsew ground input
rlabel metal3 s 0 144 800 264 6 wb_clk_i
port 2 nsew signal input
rlabel metal3 s 0 552 800 672 6 wb_rst_i
port 3 nsew signal input
rlabel metal3 s 11200 43800 12000 43920 6 wbs_hr_ack_i
port 4 nsew signal input
rlabel metal3 s 11200 1640 12000 1760 6 wbs_hr_cyc_o
port 5 nsew signal tristate
rlabel metal3 s 11200 44888 12000 45008 6 wbs_hr_dat_i[0]
port 6 nsew signal input
rlabel metal3 s 11200 56040 12000 56160 6 wbs_hr_dat_i[10]
port 7 nsew signal input
rlabel metal3 s 11200 57128 12000 57248 6 wbs_hr_dat_i[11]
port 8 nsew signal input
rlabel metal3 s 11200 58216 12000 58336 6 wbs_hr_dat_i[12]
port 9 nsew signal input
rlabel metal3 s 11200 59304 12000 59424 6 wbs_hr_dat_i[13]
port 10 nsew signal input
rlabel metal3 s 11200 60528 12000 60648 6 wbs_hr_dat_i[14]
port 11 nsew signal input
rlabel metal3 s 11200 61616 12000 61736 6 wbs_hr_dat_i[15]
port 12 nsew signal input
rlabel metal3 s 11200 62704 12000 62824 6 wbs_hr_dat_i[16]
port 13 nsew signal input
rlabel metal3 s 11200 63792 12000 63912 6 wbs_hr_dat_i[17]
port 14 nsew signal input
rlabel metal3 s 11200 64880 12000 65000 6 wbs_hr_dat_i[18]
port 15 nsew signal input
rlabel metal3 s 11200 65968 12000 66088 6 wbs_hr_dat_i[19]
port 16 nsew signal input
rlabel metal3 s 11200 45976 12000 46096 6 wbs_hr_dat_i[1]
port 17 nsew signal input
rlabel metal3 s 11200 67192 12000 67312 6 wbs_hr_dat_i[20]
port 18 nsew signal input
rlabel metal3 s 11200 68280 12000 68400 6 wbs_hr_dat_i[21]
port 19 nsew signal input
rlabel metal3 s 11200 69368 12000 69488 6 wbs_hr_dat_i[22]
port 20 nsew signal input
rlabel metal3 s 11200 70456 12000 70576 6 wbs_hr_dat_i[23]
port 21 nsew signal input
rlabel metal3 s 11200 71544 12000 71664 6 wbs_hr_dat_i[24]
port 22 nsew signal input
rlabel metal3 s 11200 72632 12000 72752 6 wbs_hr_dat_i[25]
port 23 nsew signal input
rlabel metal3 s 11200 73856 12000 73976 6 wbs_hr_dat_i[26]
port 24 nsew signal input
rlabel metal3 s 11200 74944 12000 75064 6 wbs_hr_dat_i[27]
port 25 nsew signal input
rlabel metal3 s 11200 76032 12000 76152 6 wbs_hr_dat_i[28]
port 26 nsew signal input
rlabel metal3 s 11200 77120 12000 77240 6 wbs_hr_dat_i[29]
port 27 nsew signal input
rlabel metal3 s 11200 47200 12000 47320 6 wbs_hr_dat_i[2]
port 28 nsew signal input
rlabel metal3 s 11200 78208 12000 78328 6 wbs_hr_dat_i[30]
port 29 nsew signal input
rlabel metal3 s 11200 79296 12000 79416 6 wbs_hr_dat_i[31]
port 30 nsew signal input
rlabel metal3 s 11200 48288 12000 48408 6 wbs_hr_dat_i[3]
port 31 nsew signal input
rlabel metal3 s 11200 49376 12000 49496 6 wbs_hr_dat_i[4]
port 32 nsew signal input
rlabel metal3 s 11200 50464 12000 50584 6 wbs_hr_dat_i[5]
port 33 nsew signal input
rlabel metal3 s 11200 51552 12000 51672 6 wbs_hr_dat_i[6]
port 34 nsew signal input
rlabel metal3 s 11200 52640 12000 52760 6 wbs_hr_dat_i[7]
port 35 nsew signal input
rlabel metal3 s 11200 53864 12000 53984 6 wbs_hr_dat_i[8]
port 36 nsew signal input
rlabel metal3 s 11200 54952 12000 55072 6 wbs_hr_dat_i[9]
port 37 nsew signal input
rlabel metal3 s 11200 8304 12000 8424 6 wbs_hr_dat_o[0]
port 38 nsew signal tristate
rlabel metal3 s 11200 19320 12000 19440 6 wbs_hr_dat_o[10]
port 39 nsew signal tristate
rlabel metal3 s 11200 20544 12000 20664 6 wbs_hr_dat_o[11]
port 40 nsew signal tristate
rlabel metal3 s 11200 21632 12000 21752 6 wbs_hr_dat_o[12]
port 41 nsew signal tristate
rlabel metal3 s 11200 22720 12000 22840 6 wbs_hr_dat_o[13]
port 42 nsew signal tristate
rlabel metal3 s 11200 23808 12000 23928 6 wbs_hr_dat_o[14]
port 43 nsew signal tristate
rlabel metal3 s 11200 24896 12000 25016 6 wbs_hr_dat_o[15]
port 44 nsew signal tristate
rlabel metal3 s 11200 25984 12000 26104 6 wbs_hr_dat_o[16]
port 45 nsew signal tristate
rlabel metal3 s 11200 27208 12000 27328 6 wbs_hr_dat_o[17]
port 46 nsew signal tristate
rlabel metal3 s 11200 28296 12000 28416 6 wbs_hr_dat_o[18]
port 47 nsew signal tristate
rlabel metal3 s 11200 29384 12000 29504 6 wbs_hr_dat_o[19]
port 48 nsew signal tristate
rlabel metal3 s 11200 9392 12000 9512 6 wbs_hr_dat_o[1]
port 49 nsew signal tristate
rlabel metal3 s 11200 30472 12000 30592 6 wbs_hr_dat_o[20]
port 50 nsew signal tristate
rlabel metal3 s 11200 31560 12000 31680 6 wbs_hr_dat_o[21]
port 51 nsew signal tristate
rlabel metal3 s 11200 32648 12000 32768 6 wbs_hr_dat_o[22]
port 52 nsew signal tristate
rlabel metal3 s 11200 33872 12000 33992 6 wbs_hr_dat_o[23]
port 53 nsew signal tristate
rlabel metal3 s 11200 34960 12000 35080 6 wbs_hr_dat_o[24]
port 54 nsew signal tristate
rlabel metal3 s 11200 36048 12000 36168 6 wbs_hr_dat_o[25]
port 55 nsew signal tristate
rlabel metal3 s 11200 37136 12000 37256 6 wbs_hr_dat_o[26]
port 56 nsew signal tristate
rlabel metal3 s 11200 38224 12000 38344 6 wbs_hr_dat_o[27]
port 57 nsew signal tristate
rlabel metal3 s 11200 39312 12000 39432 6 wbs_hr_dat_o[28]
port 58 nsew signal tristate
rlabel metal3 s 11200 40536 12000 40656 6 wbs_hr_dat_o[29]
port 59 nsew signal tristate
rlabel metal3 s 11200 10480 12000 10600 6 wbs_hr_dat_o[2]
port 60 nsew signal tristate
rlabel metal3 s 11200 41624 12000 41744 6 wbs_hr_dat_o[30]
port 61 nsew signal tristate
rlabel metal3 s 11200 42712 12000 42832 6 wbs_hr_dat_o[31]
port 62 nsew signal tristate
rlabel metal3 s 11200 11568 12000 11688 6 wbs_hr_dat_o[3]
port 63 nsew signal tristate
rlabel metal3 s 11200 12656 12000 12776 6 wbs_hr_dat_o[4]
port 64 nsew signal tristate
rlabel metal3 s 11200 13880 12000 14000 6 wbs_hr_dat_o[5]
port 65 nsew signal tristate
rlabel metal3 s 11200 14968 12000 15088 6 wbs_hr_dat_o[6]
port 66 nsew signal tristate
rlabel metal3 s 11200 16056 12000 16176 6 wbs_hr_dat_o[7]
port 67 nsew signal tristate
rlabel metal3 s 11200 17144 12000 17264 6 wbs_hr_dat_o[8]
port 68 nsew signal tristate
rlabel metal3 s 11200 18232 12000 18352 6 wbs_hr_dat_o[9]
port 69 nsew signal tristate
rlabel metal3 s 11200 3816 12000 3936 6 wbs_hr_sel_o[0]
port 70 nsew signal tristate
rlabel metal3 s 11200 4904 12000 5024 6 wbs_hr_sel_o[1]
port 71 nsew signal tristate
rlabel metal3 s 11200 5992 12000 6112 6 wbs_hr_sel_o[2]
port 72 nsew signal tristate
rlabel metal3 s 11200 7216 12000 7336 6 wbs_hr_sel_o[3]
port 73 nsew signal tristate
rlabel metal3 s 11200 552 12000 672 6 wbs_hr_stb_o
port 74 nsew signal tristate
rlabel metal3 s 11200 2728 12000 2848 6 wbs_hr_we_o
port 75 nsew signal tristate
rlabel metal3 s 0 65152 800 65272 6 wbs_or_ack_i
port 76 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 wbs_or_cyc_o
port 77 nsew signal tristate
rlabel metal3 s 0 65696 800 65816 6 wbs_or_dat_i[0]
port 78 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 wbs_or_dat_i[10]
port 79 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 wbs_or_dat_i[11]
port 80 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 wbs_or_dat_i[12]
port 81 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 wbs_or_dat_i[13]
port 82 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 wbs_or_dat_i[14]
port 83 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 wbs_or_dat_i[15]
port 84 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 wbs_or_dat_i[16]
port 85 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 wbs_or_dat_i[17]
port 86 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 wbs_or_dat_i[18]
port 87 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 wbs_or_dat_i[19]
port 88 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 wbs_or_dat_i[1]
port 89 nsew signal input
rlabel metal3 s 0 74672 800 74792 6 wbs_or_dat_i[20]
port 90 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 wbs_or_dat_i[21]
port 91 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 wbs_or_dat_i[22]
port 92 nsew signal input
rlabel metal3 s 0 76032 800 76152 6 wbs_or_dat_i[23]
port 93 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 wbs_or_dat_i[24]
port 94 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 wbs_or_dat_i[25]
port 95 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 wbs_or_dat_i[26]
port 96 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 wbs_or_dat_i[27]
port 97 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 wbs_or_dat_i[28]
port 98 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 wbs_or_dat_i[29]
port 99 nsew signal input
rlabel metal3 s 0 66512 800 66632 6 wbs_or_dat_i[2]
port 100 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 wbs_or_dat_i[30]
port 101 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 wbs_or_dat_i[31]
port 102 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 wbs_or_dat_i[3]
port 103 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 wbs_or_dat_i[4]
port 104 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 wbs_or_dat_i[5]
port 105 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 wbs_or_dat_i[6]
port 106 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 wbs_or_dat_i[7]
port 107 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 wbs_or_dat_i[8]
port 108 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 wbs_or_dat_i[9]
port 109 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 wbs_or_dat_o[0]
port 110 nsew signal tristate
rlabel metal3 s 0 55360 800 55480 6 wbs_or_dat_o[10]
port 111 nsew signal tristate
rlabel metal3 s 0 55768 800 55888 6 wbs_or_dat_o[11]
port 112 nsew signal tristate
rlabel metal3 s 0 56176 800 56296 6 wbs_or_dat_o[12]
port 113 nsew signal tristate
rlabel metal3 s 0 56720 800 56840 6 wbs_or_dat_o[13]
port 114 nsew signal tristate
rlabel metal3 s 0 57128 800 57248 6 wbs_or_dat_o[14]
port 115 nsew signal tristate
rlabel metal3 s 0 57536 800 57656 6 wbs_or_dat_o[15]
port 116 nsew signal tristate
rlabel metal3 s 0 58080 800 58200 6 wbs_or_dat_o[16]
port 117 nsew signal tristate
rlabel metal3 s 0 58488 800 58608 6 wbs_or_dat_o[17]
port 118 nsew signal tristate
rlabel metal3 s 0 58896 800 59016 6 wbs_or_dat_o[18]
port 119 nsew signal tristate
rlabel metal3 s 0 59440 800 59560 6 wbs_or_dat_o[19]
port 120 nsew signal tristate
rlabel metal3 s 0 51280 800 51400 6 wbs_or_dat_o[1]
port 121 nsew signal tristate
rlabel metal3 s 0 59848 800 59968 6 wbs_or_dat_o[20]
port 122 nsew signal tristate
rlabel metal3 s 0 60256 800 60376 6 wbs_or_dat_o[21]
port 123 nsew signal tristate
rlabel metal3 s 0 60664 800 60784 6 wbs_or_dat_o[22]
port 124 nsew signal tristate
rlabel metal3 s 0 61208 800 61328 6 wbs_or_dat_o[23]
port 125 nsew signal tristate
rlabel metal3 s 0 61616 800 61736 6 wbs_or_dat_o[24]
port 126 nsew signal tristate
rlabel metal3 s 0 62024 800 62144 6 wbs_or_dat_o[25]
port 127 nsew signal tristate
rlabel metal3 s 0 62568 800 62688 6 wbs_or_dat_o[26]
port 128 nsew signal tristate
rlabel metal3 s 0 62976 800 63096 6 wbs_or_dat_o[27]
port 129 nsew signal tristate
rlabel metal3 s 0 63384 800 63504 6 wbs_or_dat_o[28]
port 130 nsew signal tristate
rlabel metal3 s 0 63928 800 64048 6 wbs_or_dat_o[29]
port 131 nsew signal tristate
rlabel metal3 s 0 51688 800 51808 6 wbs_or_dat_o[2]
port 132 nsew signal tristate
rlabel metal3 s 0 64336 800 64456 6 wbs_or_dat_o[30]
port 133 nsew signal tristate
rlabel metal3 s 0 64744 800 64864 6 wbs_or_dat_o[31]
port 134 nsew signal tristate
rlabel metal3 s 0 52232 800 52352 6 wbs_or_dat_o[3]
port 135 nsew signal tristate
rlabel metal3 s 0 52640 800 52760 6 wbs_or_dat_o[4]
port 136 nsew signal tristate
rlabel metal3 s 0 53048 800 53168 6 wbs_or_dat_o[5]
port 137 nsew signal tristate
rlabel metal3 s 0 53592 800 53712 6 wbs_or_dat_o[6]
port 138 nsew signal tristate
rlabel metal3 s 0 54000 800 54120 6 wbs_or_dat_o[7]
port 139 nsew signal tristate
rlabel metal3 s 0 54408 800 54528 6 wbs_or_dat_o[8]
port 140 nsew signal tristate
rlabel metal3 s 0 54952 800 55072 6 wbs_or_dat_o[9]
port 141 nsew signal tristate
rlabel metal3 s 0 49104 800 49224 6 wbs_or_sel_o[0]
port 142 nsew signal tristate
rlabel metal3 s 0 49512 800 49632 6 wbs_or_sel_o[1]
port 143 nsew signal tristate
rlabel metal3 s 0 49920 800 50040 6 wbs_or_sel_o[2]
port 144 nsew signal tristate
rlabel metal3 s 0 50328 800 50448 6 wbs_or_sel_o[3]
port 145 nsew signal tristate
rlabel metal3 s 0 47744 800 47864 6 wbs_or_stb_o
port 146 nsew signal tristate
rlabel metal3 s 0 48560 800 48680 6 wbs_or_we_o
port 147 nsew signal tristate
rlabel metal3 s 0 32920 800 33040 6 wbs_ufp_ack_o
port 148 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 wbs_ufp_adr_i[0]
port 149 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 wbs_ufp_adr_i[10]
port 150 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 wbs_ufp_adr_i[11]
port 151 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wbs_ufp_adr_i[12]
port 152 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 wbs_ufp_adr_i[13]
port 153 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 wbs_ufp_adr_i[14]
port 154 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wbs_ufp_adr_i[15]
port 155 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 wbs_ufp_adr_i[16]
port 156 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 wbs_ufp_adr_i[17]
port 157 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 wbs_ufp_adr_i[18]
port 158 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 wbs_ufp_adr_i[19]
port 159 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 wbs_ufp_adr_i[1]
port 160 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 wbs_ufp_adr_i[20]
port 161 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 wbs_ufp_adr_i[21]
port 162 nsew signal input
rlabel metal3 s 0 14016 800 14136 6 wbs_ufp_adr_i[22]
port 163 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 wbs_ufp_adr_i[23]
port 164 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 wbs_ufp_adr_i[24]
port 165 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 wbs_ufp_adr_i[25]
port 166 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wbs_ufp_adr_i[26]
port 167 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 wbs_ufp_adr_i[27]
port 168 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 wbs_ufp_adr_i[28]
port 169 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 wbs_ufp_adr_i[29]
port 170 nsew signal input
rlabel metal3 s 0 5040 800 5160 6 wbs_ufp_adr_i[2]
port 171 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 wbs_ufp_adr_i[30]
port 172 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wbs_ufp_adr_i[31]
port 173 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 wbs_ufp_adr_i[3]
port 174 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 wbs_ufp_adr_i[4]
port 175 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 wbs_ufp_adr_i[5]
port 176 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wbs_ufp_adr_i[6]
port 177 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 wbs_ufp_adr_i[7]
port 178 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 wbs_ufp_adr_i[8]
port 179 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 wbs_ufp_adr_i[9]
port 180 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 wbs_ufp_cyc_i
port 181 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 wbs_ufp_dat_i[0]
port 182 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 wbs_ufp_dat_i[10]
port 183 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 wbs_ufp_dat_i[11]
port 184 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 wbs_ufp_dat_i[12]
port 185 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 wbs_ufp_dat_i[13]
port 186 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 wbs_ufp_dat_i[14]
port 187 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wbs_ufp_dat_i[15]
port 188 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wbs_ufp_dat_i[16]
port 189 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 wbs_ufp_dat_i[17]
port 190 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wbs_ufp_dat_i[18]
port 191 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 wbs_ufp_dat_i[19]
port 192 nsew signal input
rlabel metal3 s 0 18912 800 19032 6 wbs_ufp_dat_i[1]
port 193 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 wbs_ufp_dat_i[20]
port 194 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 wbs_ufp_dat_i[21]
port 195 nsew signal input
rlabel metal3 s 0 28432 800 28552 6 wbs_ufp_dat_i[22]
port 196 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 wbs_ufp_dat_i[23]
port 197 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 wbs_ufp_dat_i[24]
port 198 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 wbs_ufp_dat_i[25]
port 199 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 wbs_ufp_dat_i[26]
port 200 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 wbs_ufp_dat_i[27]
port 201 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 wbs_ufp_dat_i[28]
port 202 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 wbs_ufp_dat_i[29]
port 203 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wbs_ufp_dat_i[2]
port 204 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 wbs_ufp_dat_i[30]
port 205 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 wbs_ufp_dat_i[31]
port 206 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 wbs_ufp_dat_i[3]
port 207 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wbs_ufp_dat_i[4]
port 208 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wbs_ufp_dat_i[5]
port 209 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 wbs_ufp_dat_i[6]
port 210 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 wbs_ufp_dat_i[7]
port 211 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 wbs_ufp_dat_i[8]
port 212 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 wbs_ufp_dat_i[9]
port 213 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 wbs_ufp_dat_o[0]
port 214 nsew signal tristate
rlabel metal3 s 0 37816 800 37936 6 wbs_ufp_dat_o[10]
port 215 nsew signal tristate
rlabel metal3 s 0 38224 800 38344 6 wbs_ufp_dat_o[11]
port 216 nsew signal tristate
rlabel metal3 s 0 38768 800 38888 6 wbs_ufp_dat_o[12]
port 217 nsew signal tristate
rlabel metal3 s 0 39176 800 39296 6 wbs_ufp_dat_o[13]
port 218 nsew signal tristate
rlabel metal3 s 0 39584 800 39704 6 wbs_ufp_dat_o[14]
port 219 nsew signal tristate
rlabel metal3 s 0 40128 800 40248 6 wbs_ufp_dat_o[15]
port 220 nsew signal tristate
rlabel metal3 s 0 40536 800 40656 6 wbs_ufp_dat_o[16]
port 221 nsew signal tristate
rlabel metal3 s 0 40944 800 41064 6 wbs_ufp_dat_o[17]
port 222 nsew signal tristate
rlabel metal3 s 0 41352 800 41472 6 wbs_ufp_dat_o[18]
port 223 nsew signal tristate
rlabel metal3 s 0 41896 800 42016 6 wbs_ufp_dat_o[19]
port 224 nsew signal tristate
rlabel metal3 s 0 33736 800 33856 6 wbs_ufp_dat_o[1]
port 225 nsew signal tristate
rlabel metal3 s 0 42304 800 42424 6 wbs_ufp_dat_o[20]
port 226 nsew signal tristate
rlabel metal3 s 0 42712 800 42832 6 wbs_ufp_dat_o[21]
port 227 nsew signal tristate
rlabel metal3 s 0 43256 800 43376 6 wbs_ufp_dat_o[22]
port 228 nsew signal tristate
rlabel metal3 s 0 43664 800 43784 6 wbs_ufp_dat_o[23]
port 229 nsew signal tristate
rlabel metal3 s 0 44072 800 44192 6 wbs_ufp_dat_o[24]
port 230 nsew signal tristate
rlabel metal3 s 0 44616 800 44736 6 wbs_ufp_dat_o[25]
port 231 nsew signal tristate
rlabel metal3 s 0 45024 800 45144 6 wbs_ufp_dat_o[26]
port 232 nsew signal tristate
rlabel metal3 s 0 45432 800 45552 6 wbs_ufp_dat_o[27]
port 233 nsew signal tristate
rlabel metal3 s 0 45840 800 45960 6 wbs_ufp_dat_o[28]
port 234 nsew signal tristate
rlabel metal3 s 0 46384 800 46504 6 wbs_ufp_dat_o[29]
port 235 nsew signal tristate
rlabel metal3 s 0 34280 800 34400 6 wbs_ufp_dat_o[2]
port 236 nsew signal tristate
rlabel metal3 s 0 46792 800 46912 6 wbs_ufp_dat_o[30]
port 237 nsew signal tristate
rlabel metal3 s 0 47200 800 47320 6 wbs_ufp_dat_o[31]
port 238 nsew signal tristate
rlabel metal3 s 0 34688 800 34808 6 wbs_ufp_dat_o[3]
port 239 nsew signal tristate
rlabel metal3 s 0 35096 800 35216 6 wbs_ufp_dat_o[4]
port 240 nsew signal tristate
rlabel metal3 s 0 35504 800 35624 6 wbs_ufp_dat_o[5]
port 241 nsew signal tristate
rlabel metal3 s 0 36048 800 36168 6 wbs_ufp_dat_o[6]
port 242 nsew signal tristate
rlabel metal3 s 0 36456 800 36576 6 wbs_ufp_dat_o[7]
port 243 nsew signal tristate
rlabel metal3 s 0 36864 800 36984 6 wbs_ufp_dat_o[8]
port 244 nsew signal tristate
rlabel metal3 s 0 37408 800 37528 6 wbs_ufp_dat_o[9]
port 245 nsew signal tristate
rlabel metal3 s 0 2320 800 2440 6 wbs_ufp_sel_i[0]
port 246 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 wbs_ufp_sel_i[1]
port 247 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 wbs_ufp_sel_i[2]
port 248 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 wbs_ufp_sel_i[3]
port 249 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wbs_ufp_stb_i
port 250 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 wbs_ufp_we_i
port 251 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12000 80000
<< end >>
