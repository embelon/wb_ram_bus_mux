magic
tech sky130A
magscale 1 2
timestamp 1636573153
<< locali >>
rect 10977 76619 11011 78625
rect 11069 73083 11103 77469
rect 9781 65943 9815 66181
rect 10885 65943 10919 66249
rect 10977 66011 11011 69377
rect 11069 66215 11103 69853
rect 10885 65909 11011 65943
rect 857 48535 891 54145
rect 949 51459 983 64617
rect 2697 62883 2731 62985
rect 2789 56695 2823 57001
rect 857 41531 891 45509
rect 949 39491 983 42313
rect 3801 40511 3835 40681
rect 10977 32011 11011 65909
rect 11069 57579 11103 60673
rect 11069 51867 11103 55709
rect 11161 51595 11195 57885
rect 11253 56491 11287 61761
rect 11253 51459 11287 56321
rect 11345 50779 11379 57409
rect 11437 55335 11471 62237
rect 11529 50439 11563 58497
rect 10977 26299 11011 28917
rect 10919 26197 11011 26231
rect 10977 22559 11011 26197
rect 10977 22151 11011 22525
rect 10977 2499 11011 5729
<< viali >>
rect 10977 78625 11011 78659
rect 9321 77673 9355 77707
rect 2697 77605 2731 77639
rect 1409 77469 1443 77503
rect 2053 77469 2087 77503
rect 2881 77469 2915 77503
rect 3801 77469 3835 77503
rect 9137 77469 9171 77503
rect 9873 77469 9907 77503
rect 1593 77333 1627 77367
rect 2237 77333 2271 77367
rect 3985 77333 4019 77367
rect 10057 77333 10091 77367
rect 9321 77129 9355 77163
rect 1409 76993 1443 77027
rect 2053 76993 2087 77027
rect 2697 76993 2731 77027
rect 9137 76993 9171 77027
rect 9873 76993 9907 77027
rect 1593 76789 1627 76823
rect 2237 76789 2271 76823
rect 2881 76789 2915 76823
rect 10057 76789 10091 76823
rect 10057 76585 10091 76619
rect 10977 76585 11011 76619
rect 11069 77469 11103 77503
rect 1409 76381 1443 76415
rect 9873 76381 9907 76415
rect 1593 76245 1627 76279
rect 1593 76041 1627 76075
rect 1409 75905 1443 75939
rect 9873 75905 9907 75939
rect 10057 75701 10091 75735
rect 1593 75429 1627 75463
rect 1409 75293 1443 75327
rect 2053 75293 2087 75327
rect 9873 75293 9907 75327
rect 2237 75157 2271 75191
rect 10057 75157 10091 75191
rect 2973 74953 3007 74987
rect 1593 74885 1627 74919
rect 1685 74885 1719 74919
rect 2697 74885 2731 74919
rect 1409 74817 1443 74851
rect 1777 74817 1811 74851
rect 2421 74817 2455 74851
rect 2605 74817 2639 74851
rect 2789 74817 2823 74851
rect 1961 74613 1995 74647
rect 1961 74409 1995 74443
rect 2973 74341 3007 74375
rect 1409 74205 1443 74239
rect 1685 74205 1719 74239
rect 1777 74205 1811 74239
rect 2421 74205 2455 74239
rect 2697 74205 2731 74239
rect 2789 74205 2823 74239
rect 3801 74205 3835 74239
rect 9873 74205 9907 74239
rect 1593 74137 1627 74171
rect 2605 74137 2639 74171
rect 3985 74069 4019 74103
rect 10057 74069 10091 74103
rect 3065 73865 3099 73899
rect 4077 73865 4111 73899
rect 5089 73865 5123 73899
rect 1685 73797 1719 73831
rect 2697 73797 2731 73831
rect 2789 73797 2823 73831
rect 3801 73797 3835 73831
rect 4721 73797 4755 73831
rect 1409 73729 1443 73763
rect 1593 73729 1627 73763
rect 1777 73729 1811 73763
rect 2513 73729 2547 73763
rect 2881 73729 2915 73763
rect 3525 73729 3559 73763
rect 3709 73729 3743 73763
rect 3893 73729 3927 73763
rect 4557 73729 4591 73763
rect 4809 73729 4843 73763
rect 4951 73729 4985 73763
rect 9873 73729 9907 73763
rect 1961 73525 1995 73559
rect 10057 73525 10091 73559
rect 3065 73253 3099 73287
rect 1409 73117 1443 73151
rect 1685 73117 1719 73151
rect 1777 73117 1811 73151
rect 2513 73117 2547 73151
rect 2881 73117 2915 73151
rect 9873 73117 9907 73151
rect 1593 73049 1627 73083
rect 2697 73049 2731 73083
rect 2789 73049 2823 73083
rect 11069 73049 11103 73083
rect 1961 72981 1995 73015
rect 10057 72981 10091 73015
rect 1409 72641 1443 72675
rect 2053 72641 2087 72675
rect 2973 72641 3007 72675
rect 4261 72641 4295 72675
rect 2697 72573 2731 72607
rect 3985 72573 4019 72607
rect 1593 72437 1627 72471
rect 2237 72437 2271 72471
rect 1593 72233 1627 72267
rect 4353 72165 4387 72199
rect 1409 72029 1443 72063
rect 2513 72029 2547 72063
rect 2697 72029 2731 72063
rect 2789 72029 2823 72063
rect 2881 72029 2915 72063
rect 3801 72029 3835 72063
rect 4077 72029 4111 72063
rect 4169 72029 4203 72063
rect 9873 72029 9907 72063
rect 3985 71961 4019 71995
rect 3065 71893 3099 71927
rect 10057 71893 10091 71927
rect 2329 71621 2363 71655
rect 1409 71553 1443 71587
rect 2053 71553 2087 71587
rect 2237 71553 2271 71587
rect 2421 71553 2455 71587
rect 3617 71553 3651 71587
rect 3893 71553 3927 71587
rect 9873 71553 9907 71587
rect 1593 71349 1627 71383
rect 2605 71349 2639 71383
rect 10057 71349 10091 71383
rect 3801 71009 3835 71043
rect 1409 70941 1443 70975
rect 4077 70941 4111 70975
rect 1593 70805 1627 70839
rect 1593 70601 1627 70635
rect 10057 70601 10091 70635
rect 1409 70465 1443 70499
rect 9873 70465 9907 70499
rect 1409 69853 1443 69887
rect 9873 69853 9907 69887
rect 11069 69853 11103 69887
rect 1593 69717 1627 69751
rect 10057 69717 10091 69751
rect 1409 69377 1443 69411
rect 9873 69377 9907 69411
rect 10977 69377 11011 69411
rect 1593 69173 1627 69207
rect 10057 69173 10091 69207
rect 1409 68765 1443 68799
rect 1593 68629 1627 68663
rect 1409 68289 1443 68323
rect 9873 68289 9907 68323
rect 10057 68153 10091 68187
rect 1593 68085 1627 68119
rect 1593 67881 1627 67915
rect 2053 67813 2087 67847
rect 1409 67677 1443 67711
rect 2237 67677 2271 67711
rect 9873 67677 9907 67711
rect 10057 67541 10091 67575
rect 1409 67201 1443 67235
rect 2237 67201 2271 67235
rect 9873 67201 9907 67235
rect 1593 66997 1627 67031
rect 2053 66997 2087 67031
rect 10057 66997 10091 67031
rect 2973 66793 3007 66827
rect 1409 66589 1443 66623
rect 2421 66589 2455 66623
rect 2697 66589 2731 66623
rect 2789 66589 2823 66623
rect 2605 66521 2639 66555
rect 1593 66453 1627 66487
rect 10885 66249 10919 66283
rect 1685 66181 1719 66215
rect 3709 66181 3743 66215
rect 9781 66181 9815 66215
rect 1409 66113 1443 66147
rect 1593 66113 1627 66147
rect 1777 66113 1811 66147
rect 2421 66113 2455 66147
rect 2559 66113 2593 66147
rect 2697 66113 2731 66147
rect 2789 66113 2823 66147
rect 3433 66113 3467 66147
rect 3617 66113 3651 66147
rect 3801 66113 3835 66147
rect 2973 65977 3007 66011
rect 3985 65977 4019 66011
rect 9873 66113 9907 66147
rect 11069 66181 11103 66215
rect 10977 65977 11011 66011
rect 1961 65909 1995 65943
rect 9781 65909 9815 65943
rect 10057 65909 10091 65943
rect 2973 65569 3007 65603
rect 3249 65569 3283 65603
rect 4077 65569 4111 65603
rect 1409 65501 1443 65535
rect 3801 65501 3835 65535
rect 9873 65501 9907 65535
rect 1593 65365 1627 65399
rect 10057 65365 10091 65399
rect 2973 65161 3007 65195
rect 2605 65093 2639 65127
rect 1409 65025 1443 65059
rect 2421 65025 2455 65059
rect 2697 65025 2731 65059
rect 2789 65025 2823 65059
rect 1593 64889 1627 64923
rect 949 64617 983 64651
rect 2513 64617 2547 64651
rect 857 54145 891 54179
rect 2053 64549 2087 64583
rect 1501 64413 1535 64447
rect 1777 64413 1811 64447
rect 1869 64413 1903 64447
rect 2697 64413 2731 64447
rect 9873 64413 9907 64447
rect 1685 64345 1719 64379
rect 10057 64277 10091 64311
rect 3065 64073 3099 64107
rect 1777 64005 1811 64039
rect 2697 64005 2731 64039
rect 1501 63937 1535 63971
rect 1685 63937 1719 63971
rect 1915 63937 1949 63971
rect 2513 63937 2547 63971
rect 2789 63937 2823 63971
rect 2881 63937 2915 63971
rect 9873 63937 9907 63971
rect 2053 63801 2087 63835
rect 10057 63733 10091 63767
rect 2145 63461 2179 63495
rect 1593 63325 1627 63359
rect 1869 63325 1903 63359
rect 1961 63325 1995 63359
rect 2789 63325 2823 63359
rect 3985 63325 4019 63359
rect 9873 63325 9907 63359
rect 1777 63257 1811 63291
rect 2605 63189 2639 63223
rect 3801 63189 3835 63223
rect 10057 63189 10091 63223
rect 2697 62985 2731 63019
rect 1869 62917 1903 62951
rect 1685 62849 1719 62883
rect 1961 62849 1995 62883
rect 2053 62849 2087 62883
rect 2697 62849 2731 62883
rect 2789 62849 2823 62883
rect 3065 62849 3099 62883
rect 2237 62645 2271 62679
rect 2973 62305 3007 62339
rect 3249 62305 3283 62339
rect 1685 62237 1719 62271
rect 9873 62237 9907 62271
rect 1501 62101 1535 62135
rect 10057 62101 10091 62135
rect 1685 61761 1719 61795
rect 2329 61761 2363 61795
rect 9873 61761 9907 61795
rect 1501 61557 1535 61591
rect 2145 61557 2179 61591
rect 10057 61557 10091 61591
rect 1685 61149 1719 61183
rect 1501 61013 1535 61047
rect 1685 60673 1719 60707
rect 9873 60673 9907 60707
rect 10057 60537 10091 60571
rect 1501 60469 1535 60503
rect 1685 60061 1719 60095
rect 9873 60061 9907 60095
rect 1501 59925 1535 59959
rect 10057 59925 10091 59959
rect 1685 59585 1719 59619
rect 9873 59585 9907 59619
rect 1501 59381 1535 59415
rect 10057 59381 10091 59415
rect 1685 58973 1719 59007
rect 1501 58837 1535 58871
rect 1685 58497 1719 58531
rect 9873 58497 9907 58531
rect 10057 58361 10091 58395
rect 1501 58293 1535 58327
rect 1409 57885 1443 57919
rect 1685 57885 1719 57919
rect 1777 57885 1811 57919
rect 2421 57885 2455 57919
rect 9873 57885 9907 57919
rect 1593 57817 1627 57851
rect 1961 57749 1995 57783
rect 2605 57749 2639 57783
rect 10057 57749 10091 57783
rect 1685 57477 1719 57511
rect 1409 57409 1443 57443
rect 1593 57409 1627 57443
rect 1777 57409 1811 57443
rect 2697 57409 2731 57443
rect 9873 57409 9907 57443
rect 1961 57273 1995 57307
rect 2513 57205 2547 57239
rect 10057 57205 10091 57239
rect 2789 57001 2823 57035
rect 3065 57001 3099 57035
rect 1961 56933 1995 56967
rect 1409 56797 1443 56831
rect 1593 56797 1627 56831
rect 1777 56797 1811 56831
rect 1685 56729 1719 56763
rect 3801 56797 3835 56831
rect 2973 56729 3007 56763
rect 2789 56661 2823 56695
rect 3985 56661 4019 56695
rect 3985 56457 4019 56491
rect 1593 56389 1627 56423
rect 1409 56321 1443 56355
rect 1685 56321 1719 56355
rect 1777 56321 1811 56355
rect 2789 56321 2823 56355
rect 3801 56321 3835 56355
rect 9873 56321 9907 56355
rect 2513 56253 2547 56287
rect 1961 56185 1995 56219
rect 10057 56117 10091 56151
rect 2237 55777 2271 55811
rect 1961 55709 1995 55743
rect 3801 55709 3835 55743
rect 9873 55709 9907 55743
rect 3985 55573 4019 55607
rect 10057 55573 10091 55607
rect 1961 55369 1995 55403
rect 1593 55301 1627 55335
rect 1409 55233 1443 55267
rect 1685 55233 1719 55267
rect 1777 55233 1811 55267
rect 2421 55233 2455 55267
rect 2605 55097 2639 55131
rect 1685 54621 1719 54655
rect 10149 54621 10183 54655
rect 1501 54485 1535 54519
rect 9965 54485 9999 54519
rect 3801 54213 3835 54247
rect 1685 54145 1719 54179
rect 2513 54145 2547 54179
rect 3985 54145 4019 54179
rect 10149 54145 10183 54179
rect 2789 54077 2823 54111
rect 1501 53941 1535 53975
rect 9965 53941 9999 53975
rect 2053 53601 2087 53635
rect 2329 53533 2363 53567
rect 6745 53533 6779 53567
rect 10149 53533 10183 53567
rect 6561 53397 6595 53431
rect 9965 53397 9999 53431
rect 2329 53193 2363 53227
rect 2973 53193 3007 53227
rect 1685 53057 1719 53091
rect 2145 53057 2179 53091
rect 2881 53057 2915 53091
rect 3065 53057 3099 53091
rect 7205 53057 7239 53091
rect 1501 52853 1535 52887
rect 7113 52853 7147 52887
rect 2421 52649 2455 52683
rect 3065 52649 3099 52683
rect 9045 52581 9079 52615
rect 1685 52445 1719 52479
rect 2421 52445 2455 52479
rect 2599 52445 2633 52479
rect 3065 52445 3099 52479
rect 3249 52445 3283 52479
rect 9137 52445 9171 52479
rect 10149 52445 10183 52479
rect 1501 52309 1535 52343
rect 9965 52309 9999 52343
rect 3249 52105 3283 52139
rect 1593 52037 1627 52071
rect 1409 51969 1443 52003
rect 1685 51969 1719 52003
rect 1777 51969 1811 52003
rect 2421 51969 2455 52003
rect 3157 51969 3191 52003
rect 3341 51969 3375 52003
rect 10149 51969 10183 52003
rect 1961 51833 1995 51867
rect 2605 51833 2639 51867
rect 9965 51765 9999 51799
rect 2973 51561 3007 51595
rect 1961 51493 1995 51527
rect 949 51425 983 51459
rect 1409 51357 1443 51391
rect 1593 51357 1627 51391
rect 1685 51357 1719 51391
rect 1823 51357 1857 51391
rect 2421 51357 2455 51391
rect 2789 51357 2823 51391
rect 4353 51357 4387 51391
rect 2605 51289 2639 51323
rect 2697 51289 2731 51323
rect 4169 51221 4203 51255
rect 3249 51017 3283 51051
rect 1685 50949 1719 50983
rect 1409 50881 1443 50915
rect 1593 50881 1627 50915
rect 1777 50881 1811 50915
rect 2421 50881 2455 50915
rect 3157 50881 3191 50915
rect 3341 50881 3375 50915
rect 4077 50881 4111 50915
rect 4721 50881 4755 50915
rect 4905 50881 4939 50915
rect 10149 50881 10183 50915
rect 2605 50745 2639 50779
rect 1961 50677 1995 50711
rect 4077 50677 4111 50711
rect 4721 50677 4755 50711
rect 9965 50677 9999 50711
rect 1961 50405 1995 50439
rect 1409 50269 1443 50303
rect 1685 50269 1719 50303
rect 1777 50269 1811 50303
rect 2697 50269 2731 50303
rect 4261 50269 4295 50303
rect 10149 50269 10183 50303
rect 1593 50201 1627 50235
rect 2513 50133 2547 50167
rect 4077 50133 4111 50167
rect 9965 50133 9999 50167
rect 2421 49929 2455 49963
rect 4077 49929 4111 49963
rect 1685 49793 1719 49827
rect 2329 49793 2363 49827
rect 2513 49793 2547 49827
rect 3433 49793 3467 49827
rect 4261 49793 4295 49827
rect 10149 49793 10183 49827
rect 1501 49657 1535 49691
rect 3249 49589 3283 49623
rect 9965 49589 9999 49623
rect 2329 49385 2363 49419
rect 3985 49249 4019 49283
rect 1685 49181 1719 49215
rect 2329 49181 2363 49215
rect 2513 49181 2547 49215
rect 4261 49181 4295 49215
rect 1501 49045 1535 49079
rect 3801 48841 3835 48875
rect 1685 48705 1719 48739
rect 3985 48705 4019 48739
rect 10149 48705 10183 48739
rect 1501 48569 1535 48603
rect 857 48501 891 48535
rect 9965 48501 9999 48535
rect 1685 48093 1719 48127
rect 10149 48093 10183 48127
rect 1501 47957 1535 47991
rect 9965 47957 9999 47991
rect 1685 47617 1719 47651
rect 3341 47617 3375 47651
rect 4353 47617 4387 47651
rect 3617 47549 3651 47583
rect 1501 47481 1535 47515
rect 4169 47413 4203 47447
rect 1501 47141 1535 47175
rect 1685 47005 1719 47039
rect 10149 47005 10183 47039
rect 9965 46869 9999 46903
rect 2237 46665 2271 46699
rect 1685 46529 1719 46563
rect 2145 46529 2179 46563
rect 2329 46529 2363 46563
rect 3709 46529 3743 46563
rect 10149 46529 10183 46563
rect 3709 46393 3743 46427
rect 1501 46325 1535 46359
rect 9965 46325 9999 46359
rect 2145 46121 2179 46155
rect 2973 46121 3007 46155
rect 1685 45917 1719 45951
rect 2145 45917 2179 45951
rect 2329 45917 2363 45951
rect 2789 45917 2823 45951
rect 2973 45917 3007 45951
rect 4077 45917 4111 45951
rect 10149 45917 10183 45951
rect 3801 45849 3835 45883
rect 1501 45781 1535 45815
rect 9965 45781 9999 45815
rect 857 45509 891 45543
rect 1685 45441 1719 45475
rect 2973 45441 3007 45475
rect 4261 45441 4295 45475
rect 2697 45373 2731 45407
rect 1501 45237 1535 45271
rect 4077 45237 4111 45271
rect 2145 45033 2179 45067
rect 2789 45033 2823 45067
rect 1685 44829 1719 44863
rect 2145 44829 2179 44863
rect 2329 44829 2363 44863
rect 2789 44829 2823 44863
rect 2973 44829 3007 44863
rect 4261 44829 4295 44863
rect 10149 44829 10183 44863
rect 3985 44761 4019 44795
rect 1501 44693 1535 44727
rect 9965 44693 9999 44727
rect 1685 44353 1719 44387
rect 10149 44353 10183 44387
rect 1501 44149 1535 44183
rect 9965 44149 9999 44183
rect 1685 43741 1719 43775
rect 10149 43741 10183 43775
rect 1501 43605 1535 43639
rect 9965 43605 9999 43639
rect 1685 43265 1719 43299
rect 3801 43265 3835 43299
rect 1501 43061 1535 43095
rect 3617 43061 3651 43095
rect 4077 42721 4111 42755
rect 1685 42653 1719 42687
rect 3801 42653 3835 42687
rect 10149 42653 10183 42687
rect 1501 42517 1535 42551
rect 9965 42517 9999 42551
rect 857 41497 891 41531
rect 949 42313 983 42347
rect 1685 42177 1719 42211
rect 3985 42177 4019 42211
rect 10149 42177 10183 42211
rect 1501 41973 1535 42007
rect 3985 41973 4019 42007
rect 9965 41973 9999 42007
rect 2145 41769 2179 41803
rect 1685 41565 1719 41599
rect 2145 41565 2179 41599
rect 2329 41565 2363 41599
rect 4077 41565 4111 41599
rect 3801 41497 3835 41531
rect 1501 41429 1535 41463
rect 2237 41225 2271 41259
rect 2881 41157 2915 41191
rect 1685 41089 1719 41123
rect 2145 41089 2179 41123
rect 2329 41089 2363 41123
rect 2789 41089 2823 41123
rect 2973 41089 3007 41123
rect 4077 41089 4111 41123
rect 10149 41089 10183 41123
rect 1501 40885 1535 40919
rect 4169 40885 4203 40919
rect 9965 40885 9999 40919
rect 2145 40681 2179 40715
rect 2789 40681 2823 40715
rect 3801 40681 3835 40715
rect 1685 40477 1719 40511
rect 2145 40477 2179 40511
rect 2329 40477 2363 40511
rect 2789 40477 2823 40511
rect 2973 40477 3007 40511
rect 3801 40477 3835 40511
rect 4077 40477 4111 40511
rect 10149 40477 10183 40511
rect 1501 40341 1535 40375
rect 3985 40341 4019 40375
rect 9965 40341 9999 40375
rect 1409 40001 1443 40035
rect 2605 40001 2639 40035
rect 2881 40001 2915 40035
rect 4169 40001 4203 40035
rect 10149 40001 10183 40035
rect 1593 39865 1627 39899
rect 3985 39797 4019 39831
rect 9965 39797 9999 39831
rect 2145 39593 2179 39627
rect 1593 39525 1627 39559
rect 949 39457 983 39491
rect 1409 39389 1443 39423
rect 2145 39389 2179 39423
rect 2329 39389 2363 39423
rect 4077 39389 4111 39423
rect 3801 39321 3835 39355
rect 1593 39049 1627 39083
rect 2237 39049 2271 39083
rect 2881 39049 2915 39083
rect 1409 38913 1443 38947
rect 2145 38913 2179 38947
rect 2329 38913 2363 38947
rect 2789 38913 2823 38947
rect 2973 38913 3007 38947
rect 10149 38913 10183 38947
rect 9965 38709 9999 38743
rect 2145 38505 2179 38539
rect 2789 38505 2823 38539
rect 1593 38437 1627 38471
rect 1409 38301 1443 38335
rect 2145 38301 2179 38335
rect 2329 38301 2363 38335
rect 2789 38301 2823 38335
rect 2973 38301 3007 38335
rect 4077 38301 4111 38335
rect 10149 38301 10183 38335
rect 3893 38165 3927 38199
rect 9965 38165 9999 38199
rect 1593 37961 1627 37995
rect 1409 37825 1443 37859
rect 2697 37825 2731 37859
rect 3985 37825 4019 37859
rect 2421 37757 2455 37791
rect 3985 37621 4019 37655
rect 3893 37349 3927 37383
rect 2421 37281 2455 37315
rect 1409 37213 1443 37247
rect 2697 37213 2731 37247
rect 4077 37213 4111 37247
rect 10149 37213 10183 37247
rect 1593 37077 1627 37111
rect 9965 37077 9999 37111
rect 2237 36873 2271 36907
rect 2881 36873 2915 36907
rect 1409 36737 1443 36771
rect 2145 36737 2179 36771
rect 2329 36737 2363 36771
rect 2789 36737 2823 36771
rect 2973 36737 3007 36771
rect 4077 36737 4111 36771
rect 4353 36737 4387 36771
rect 10149 36737 10183 36771
rect 1593 36533 1627 36567
rect 9965 36533 9999 36567
rect 1593 36329 1627 36363
rect 2789 36329 2823 36363
rect 2145 36261 2179 36295
rect 1409 36125 1443 36159
rect 2145 36125 2179 36159
rect 2329 36125 2363 36159
rect 2789 36125 2823 36159
rect 2973 36125 3007 36159
rect 4077 36125 4111 36159
rect 4353 36125 4387 36159
rect 10149 36125 10183 36159
rect 9965 35989 9999 36023
rect 2237 35785 2271 35819
rect 1409 35649 1443 35683
rect 2145 35649 2179 35683
rect 2329 35649 2363 35683
rect 4353 35649 4387 35683
rect 4077 35581 4111 35615
rect 1593 35513 1627 35547
rect 1593 35241 1627 35275
rect 1409 35037 1443 35071
rect 4353 35037 4387 35071
rect 10149 35037 10183 35071
rect 4169 34901 4203 34935
rect 9965 34901 9999 34935
rect 1593 34697 1627 34731
rect 4169 34697 4203 34731
rect 9965 34697 9999 34731
rect 1409 34561 1443 34595
rect 4353 34561 4387 34595
rect 10149 34561 10183 34595
rect 1593 34153 1627 34187
rect 1409 33949 1443 33983
rect 10149 33949 10183 33983
rect 9965 33813 9999 33847
rect 1593 33609 1627 33643
rect 1409 33473 1443 33507
rect 1593 33065 1627 33099
rect 1409 32861 1443 32895
rect 10149 32861 10183 32895
rect 9965 32725 9999 32759
rect 1593 32521 1627 32555
rect 2237 32521 2271 32555
rect 1409 32385 1443 32419
rect 2145 32385 2179 32419
rect 2329 32385 2363 32419
rect 10149 32385 10183 32419
rect 9965 32181 9999 32215
rect 11437 62237 11471 62271
rect 11253 61761 11287 61795
rect 11069 60673 11103 60707
rect 11069 57545 11103 57579
rect 11161 57885 11195 57919
rect 11069 55709 11103 55743
rect 11069 51833 11103 51867
rect 11253 56457 11287 56491
rect 11345 57409 11379 57443
rect 11161 51561 11195 51595
rect 11253 56321 11287 56355
rect 11253 51425 11287 51459
rect 11437 55301 11471 55335
rect 11529 58497 11563 58531
rect 11345 50745 11379 50779
rect 11529 50405 11563 50439
rect 2145 31977 2179 32011
rect 10977 31977 11011 32011
rect 1593 31909 1627 31943
rect 3249 31909 3283 31943
rect 1409 31773 1443 31807
rect 2145 31773 2179 31807
rect 2323 31773 2357 31807
rect 3249 31773 3283 31807
rect 1593 31433 1627 31467
rect 2237 31433 2271 31467
rect 3157 31433 3191 31467
rect 1409 31297 1443 31331
rect 2145 31297 2179 31331
rect 2329 31297 2363 31331
rect 3341 31297 3375 31331
rect 10149 31297 10183 31331
rect 9965 31093 9999 31127
rect 1593 30889 1627 30923
rect 2145 30889 2179 30923
rect 2789 30889 2823 30923
rect 1409 30685 1443 30719
rect 2145 30685 2179 30719
rect 2329 30685 2363 30719
rect 2789 30685 2823 30719
rect 2973 30685 3007 30719
rect 4077 30685 4111 30719
rect 10149 30685 10183 30719
rect 3893 30549 3927 30583
rect 9965 30549 9999 30583
rect 1409 30209 1443 30243
rect 2605 30209 2639 30243
rect 4077 30209 4111 30243
rect 10149 30209 10183 30243
rect 2881 30141 2915 30175
rect 1593 30073 1627 30107
rect 3985 30005 4019 30039
rect 9965 30005 9999 30039
rect 1593 29801 1627 29835
rect 2329 29665 2363 29699
rect 2605 29665 2639 29699
rect 1409 29597 1443 29631
rect 10149 29597 10183 29631
rect 9965 29461 9999 29495
rect 1593 29257 1627 29291
rect 2237 29257 2271 29291
rect 1409 29121 1443 29155
rect 2145 29121 2179 29155
rect 2329 29121 2363 29155
rect 9505 29121 9539 29155
rect 9597 29121 9631 29155
rect 9965 29121 9999 29155
rect 9873 28917 9907 28951
rect 10149 28917 10183 28951
rect 10977 28917 11011 28951
rect 2145 28713 2179 28747
rect 2789 28713 2823 28747
rect 9965 28713 9999 28747
rect 1593 28645 1627 28679
rect 1409 28509 1443 28543
rect 2151 28509 2185 28543
rect 2329 28509 2363 28543
rect 2789 28509 2823 28543
rect 2973 28509 3007 28543
rect 10149 28509 10183 28543
rect 1593 28169 1627 28203
rect 2881 28169 2915 28203
rect 1409 28033 1443 28067
rect 2145 28033 2179 28067
rect 2329 28033 2363 28067
rect 2789 28033 2823 28067
rect 2973 28033 3007 28067
rect 10149 28033 10183 28067
rect 2145 27897 2179 27931
rect 9965 27829 9999 27863
rect 1869 27625 1903 27659
rect 10149 27421 10183 27455
rect 1961 27353 1995 27387
rect 9965 27285 9999 27319
rect 10149 26945 10183 26979
rect 9965 26741 9999 26775
rect 1869 26537 1903 26571
rect 9873 26537 9907 26571
rect 10057 26401 10091 26435
rect 9873 26333 9907 26367
rect 1961 26265 1995 26299
rect 10149 26265 10183 26299
rect 10977 26265 11011 26299
rect 9689 26197 9723 26231
rect 10885 26197 10919 26231
rect 1869 25993 1903 26027
rect 10149 25993 10183 26027
rect 9781 25925 9815 25959
rect 9965 25925 9999 25959
rect 1961 25857 1995 25891
rect 1869 25449 1903 25483
rect 10149 25245 10183 25279
rect 1961 25177 1995 25211
rect 9965 25109 9999 25143
rect 1961 24769 1995 24803
rect 2513 24769 2547 24803
rect 2697 24769 2731 24803
rect 3157 24769 3191 24803
rect 3341 24769 3375 24803
rect 10149 24769 10183 24803
rect 1777 24633 1811 24667
rect 2513 24565 2547 24599
rect 3157 24565 3191 24599
rect 9965 24565 9999 24599
rect 1869 24361 1903 24395
rect 2513 24157 2547 24191
rect 2697 24157 2731 24191
rect 10149 24157 10183 24191
rect 1961 24089 1995 24123
rect 2605 24021 2639 24055
rect 9965 24021 9999 24055
rect 2053 23749 2087 23783
rect 1869 23681 1903 23715
rect 2789 23681 2823 23715
rect 2973 23681 3007 23715
rect 3433 23681 3467 23715
rect 3617 23681 3651 23715
rect 9965 23681 9999 23715
rect 2789 23545 2823 23579
rect 3433 23477 3467 23511
rect 10057 23477 10091 23511
rect 1869 23273 1903 23307
rect 9873 23273 9907 23307
rect 9781 23137 9815 23171
rect 9965 23137 9999 23171
rect 2513 23069 2547 23103
rect 2697 23069 2731 23103
rect 3801 23069 3835 23103
rect 3985 23069 4019 23103
rect 9137 23069 9171 23103
rect 1961 23001 1995 23035
rect 10149 23001 10183 23035
rect 2605 22933 2639 22967
rect 3893 22933 3927 22967
rect 9321 22933 9355 22967
rect 10057 22933 10091 22967
rect 1869 22729 1903 22763
rect 9689 22729 9723 22763
rect 1961 22593 1995 22627
rect 2697 22593 2731 22627
rect 8861 22593 8895 22627
rect 9965 22593 9999 22627
rect 10149 22593 10183 22627
rect 2973 22525 3007 22559
rect 9597 22525 9631 22559
rect 10977 22525 11011 22559
rect 9045 22389 9079 22423
rect 10977 22117 11011 22151
rect 1777 22049 1811 22083
rect 9505 22049 9539 22083
rect 1961 21981 1995 22015
rect 2519 21981 2553 22015
rect 2691 21981 2725 22015
rect 3985 21981 4019 22015
rect 9873 21981 9907 22015
rect 10057 21981 10091 22015
rect 10149 21981 10183 22015
rect 2605 21845 2639 21879
rect 3893 21845 3927 21879
rect 10149 21641 10183 21675
rect 3249 21573 3283 21607
rect 3985 21573 4019 21607
rect 1685 21505 1719 21539
rect 8953 21505 8987 21539
rect 9597 21505 9631 21539
rect 9965 21505 9999 21539
rect 1501 21369 1535 21403
rect 3157 21301 3191 21335
rect 3893 21301 3927 21335
rect 9137 21301 9171 21335
rect 9873 21301 9907 21335
rect 9229 21097 9263 21131
rect 9689 21097 9723 21131
rect 10149 21097 10183 21131
rect 9781 20961 9815 20995
rect 1685 20893 1719 20927
rect 9045 20893 9079 20927
rect 9689 20893 9723 20927
rect 9965 20893 9999 20927
rect 1501 20757 1535 20791
rect 10149 20553 10183 20587
rect 9781 20485 9815 20519
rect 1685 20417 1719 20451
rect 9965 20417 9999 20451
rect 1501 20281 1535 20315
rect 9965 20009 9999 20043
rect 1685 19805 1719 19839
rect 10149 19805 10183 19839
rect 1501 19669 1535 19703
rect 9965 19465 9999 19499
rect 1685 19329 1719 19363
rect 10149 19329 10183 19363
rect 1501 19125 1535 19159
rect 1685 18717 1719 18751
rect 1501 18581 1535 18615
rect 1685 18241 1719 18275
rect 2145 18241 2179 18275
rect 2329 18241 2363 18275
rect 1501 18037 1535 18071
rect 2145 18037 2179 18071
rect 1685 17629 1719 17663
rect 2145 17629 2179 17663
rect 2329 17629 2363 17663
rect 1501 17493 1535 17527
rect 2237 17493 2271 17527
rect 1685 17153 1719 17187
rect 2145 17153 2179 17187
rect 2329 17153 2363 17187
rect 1501 16949 1535 16983
rect 2145 16949 2179 16983
rect 2145 16677 2179 16711
rect 1685 16541 1719 16575
rect 2145 16541 2179 16575
rect 2329 16541 2363 16575
rect 2789 16541 2823 16575
rect 2973 16541 3007 16575
rect 1501 16405 1535 16439
rect 2881 16405 2915 16439
rect 1685 16065 1719 16099
rect 2145 16065 2179 16099
rect 2329 16065 2363 16099
rect 2789 16065 2823 16099
rect 2973 16065 3007 16099
rect 1501 15861 1535 15895
rect 2145 15861 2179 15895
rect 2789 15861 2823 15895
rect 1685 15453 1719 15487
rect 2145 15453 2179 15487
rect 2329 15453 2363 15487
rect 2789 15453 2823 15487
rect 2973 15453 3007 15487
rect 1501 15317 1535 15351
rect 2237 15317 2271 15351
rect 2881 15317 2915 15351
rect 1685 14977 1719 15011
rect 2145 14977 2179 15011
rect 2329 14977 2363 15011
rect 2789 14977 2823 15011
rect 2973 14977 3007 15011
rect 3433 14977 3467 15011
rect 3617 14977 3651 15011
rect 1501 14773 1535 14807
rect 2145 14773 2179 14807
rect 2789 14773 2823 14807
rect 3433 14773 3467 14807
rect 1685 14365 1719 14399
rect 2145 14365 2179 14399
rect 2329 14365 2363 14399
rect 2789 14365 2823 14399
rect 2973 14365 3007 14399
rect 3801 14365 3835 14399
rect 3985 14365 4019 14399
rect 1501 14229 1535 14263
rect 2237 14229 2271 14263
rect 2881 14229 2915 14263
rect 3893 14229 3927 14263
rect 1685 13889 1719 13923
rect 3249 13821 3283 13855
rect 3525 13821 3559 13855
rect 1501 13685 1535 13719
rect 2651 13481 2685 13515
rect 2421 13345 2455 13379
rect 1685 13277 1719 13311
rect 1501 13141 1535 13175
rect 1685 12801 1719 12835
rect 2697 12801 2731 12835
rect 2973 12801 3007 12835
rect 1501 12597 1535 12631
rect 1685 12189 1719 12223
rect 1501 12053 1535 12087
rect 1685 11713 1719 11747
rect 1501 11509 1535 11543
rect 1685 11101 1719 11135
rect 1501 10965 1535 10999
rect 1685 10625 1719 10659
rect 1501 10421 1535 10455
rect 3249 10081 3283 10115
rect 1685 10013 1719 10047
rect 2973 10013 3007 10047
rect 1501 9877 1535 9911
rect 1685 9537 1719 9571
rect 2145 9537 2179 9571
rect 1501 9333 1535 9367
rect 2329 9333 2363 9367
rect 2973 9129 3007 9163
rect 1685 8925 1719 8959
rect 2329 8925 2363 8959
rect 2513 8925 2547 8959
rect 2973 8925 3007 8959
rect 3157 8925 3191 8959
rect 1501 8789 1535 8823
rect 2421 8789 2455 8823
rect 3525 8585 3559 8619
rect 1685 8449 1719 8483
rect 2145 8449 2179 8483
rect 2329 8449 2363 8483
rect 2789 8449 2823 8483
rect 2973 8449 3007 8483
rect 3433 8449 3467 8483
rect 3617 8449 3651 8483
rect 1501 8313 1535 8347
rect 2145 8313 2179 8347
rect 2789 8245 2823 8279
rect 1685 7837 1719 7871
rect 2145 7837 2179 7871
rect 2329 7837 2363 7871
rect 2789 7837 2823 7871
rect 2973 7837 3007 7871
rect 3801 7837 3835 7871
rect 3985 7837 4019 7871
rect 1501 7701 1535 7735
rect 2237 7701 2271 7735
rect 2881 7701 2915 7735
rect 3893 7701 3927 7735
rect 1869 7497 1903 7531
rect 1961 7361 1995 7395
rect 2789 7361 2823 7395
rect 3249 7361 3283 7395
rect 3433 7361 3467 7395
rect 2605 7157 2639 7191
rect 3249 7157 3283 7191
rect 3157 6817 3191 6851
rect 1685 6749 1719 6783
rect 2881 6749 2915 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 10149 6749 10183 6783
rect 1501 6613 1535 6647
rect 3893 6613 3927 6647
rect 9965 6613 9999 6647
rect 2053 6409 2087 6443
rect 2237 6273 2271 6307
rect 2697 6273 2731 6307
rect 4261 6273 4295 6307
rect 2973 6205 3007 6239
rect 4077 6137 4111 6171
rect 3249 5865 3283 5899
rect 4721 5865 4755 5899
rect 3893 5729 3927 5763
rect 10977 5729 11011 5763
rect 1685 5661 1719 5695
rect 2145 5661 2179 5695
rect 2329 5661 2363 5695
rect 3249 5661 3283 5695
rect 4077 5661 4111 5695
rect 4905 5661 4939 5695
rect 10149 5661 10183 5695
rect 1501 5525 1535 5559
rect 2237 5525 2271 5559
rect 9965 5525 9999 5559
rect 9965 5321 9999 5355
rect 1685 5185 1719 5219
rect 2145 5185 2179 5219
rect 2329 5185 2363 5219
rect 2789 5185 2823 5219
rect 2973 5185 3007 5219
rect 3893 5185 3927 5219
rect 4077 5185 4111 5219
rect 10149 5185 10183 5219
rect 2145 5049 2179 5083
rect 1501 4981 1535 5015
rect 2789 4981 2823 5015
rect 1685 4573 1719 4607
rect 2145 4573 2179 4607
rect 2329 4573 2363 4607
rect 2789 4573 2823 4607
rect 2973 4573 3007 4607
rect 1501 4437 1535 4471
rect 2237 4437 2271 4471
rect 2881 4437 2915 4471
rect 9965 4233 9999 4267
rect 1685 4097 1719 4131
rect 2145 4097 2179 4131
rect 10149 4097 10183 4131
rect 1501 3893 1535 3927
rect 2329 3893 2363 3927
rect 9965 3689 9999 3723
rect 1685 3485 1719 3519
rect 2329 3485 2363 3519
rect 10149 3485 10183 3519
rect 1501 3349 1535 3383
rect 2145 3349 2179 3383
rect 1685 3009 1719 3043
rect 9873 3009 9907 3043
rect 10149 2941 10183 2975
rect 1501 2805 1535 2839
rect 9873 2465 9907 2499
rect 10977 2465 11011 2499
rect 1685 2397 1719 2431
rect 2145 2397 2179 2431
rect 2881 2397 2915 2431
rect 10149 2397 10183 2431
rect 1501 2261 1535 2295
rect 2329 2261 2363 2295
rect 3065 2261 3099 2295
<< metal1 >>
rect 10962 78656 10968 78668
rect 10923 78628 10968 78656
rect 10962 78616 10968 78628
rect 11020 78616 11026 78668
rect 1104 77818 10856 77840
rect 1104 77766 2582 77818
rect 2634 77766 2646 77818
rect 2698 77766 2710 77818
rect 2762 77766 2774 77818
rect 2826 77766 2838 77818
rect 2890 77766 5845 77818
rect 5897 77766 5909 77818
rect 5961 77766 5973 77818
rect 6025 77766 6037 77818
rect 6089 77766 6101 77818
rect 6153 77766 9109 77818
rect 9161 77766 9173 77818
rect 9225 77766 9237 77818
rect 9289 77766 9301 77818
rect 9353 77766 9365 77818
rect 9417 77766 10856 77818
rect 1104 77744 10856 77766
rect 9309 77707 9367 77713
rect 9309 77673 9321 77707
rect 9355 77704 9367 77707
rect 9490 77704 9496 77716
rect 9355 77676 9496 77704
rect 9355 77673 9367 77676
rect 9309 77667 9367 77673
rect 9490 77664 9496 77676
rect 9548 77664 9554 77716
rect 1762 77596 1768 77648
rect 1820 77636 1826 77648
rect 2685 77639 2743 77645
rect 2685 77636 2697 77639
rect 1820 77608 2697 77636
rect 1820 77596 1826 77608
rect 2685 77605 2697 77608
rect 2731 77605 2743 77639
rect 2685 77599 2743 77605
rect 1394 77500 1400 77512
rect 1355 77472 1400 77500
rect 1394 77460 1400 77472
rect 1452 77460 1458 77512
rect 2038 77500 2044 77512
rect 1999 77472 2044 77500
rect 2038 77460 2044 77472
rect 2096 77460 2102 77512
rect 2869 77503 2927 77509
rect 2869 77469 2881 77503
rect 2915 77500 2927 77503
rect 2958 77500 2964 77512
rect 2915 77472 2964 77500
rect 2915 77469 2927 77472
rect 2869 77463 2927 77469
rect 2958 77460 2964 77472
rect 3016 77460 3022 77512
rect 3786 77500 3792 77512
rect 3747 77472 3792 77500
rect 3786 77460 3792 77472
rect 3844 77460 3850 77512
rect 5534 77460 5540 77512
rect 5592 77500 5598 77512
rect 9125 77503 9183 77509
rect 9125 77500 9137 77503
rect 5592 77472 9137 77500
rect 5592 77460 5598 77472
rect 9125 77469 9137 77472
rect 9171 77469 9183 77503
rect 9125 77463 9183 77469
rect 9861 77503 9919 77509
rect 9861 77469 9873 77503
rect 9907 77500 9919 77503
rect 11057 77503 11115 77509
rect 11057 77500 11069 77503
rect 9907 77472 11069 77500
rect 9907 77469 9919 77472
rect 9861 77463 9919 77469
rect 11057 77469 11069 77472
rect 11103 77469 11115 77503
rect 11057 77463 11115 77469
rect 1581 77367 1639 77373
rect 1581 77333 1593 77367
rect 1627 77364 1639 77367
rect 1670 77364 1676 77376
rect 1627 77336 1676 77364
rect 1627 77333 1639 77336
rect 1581 77327 1639 77333
rect 1670 77324 1676 77336
rect 1728 77324 1734 77376
rect 2225 77367 2283 77373
rect 2225 77333 2237 77367
rect 2271 77364 2283 77367
rect 2498 77364 2504 77376
rect 2271 77336 2504 77364
rect 2271 77333 2283 77336
rect 2225 77327 2283 77333
rect 2498 77324 2504 77336
rect 2556 77324 2562 77376
rect 3970 77364 3976 77376
rect 3931 77336 3976 77364
rect 3970 77324 3976 77336
rect 4028 77324 4034 77376
rect 10042 77364 10048 77376
rect 10003 77336 10048 77364
rect 10042 77324 10048 77336
rect 10100 77324 10106 77376
rect 1104 77274 10856 77296
rect 1104 77222 4213 77274
rect 4265 77222 4277 77274
rect 4329 77222 4341 77274
rect 4393 77222 4405 77274
rect 4457 77222 4469 77274
rect 4521 77222 7477 77274
rect 7529 77222 7541 77274
rect 7593 77222 7605 77274
rect 7657 77222 7669 77274
rect 7721 77222 7733 77274
rect 7785 77222 10856 77274
rect 1104 77200 10856 77222
rect 9309 77163 9367 77169
rect 9309 77129 9321 77163
rect 9355 77160 9367 77163
rect 9582 77160 9588 77172
rect 9355 77132 9588 77160
rect 9355 77129 9367 77132
rect 9309 77123 9367 77129
rect 9582 77120 9588 77132
rect 9640 77120 9646 77172
rect 1302 76984 1308 77036
rect 1360 77024 1366 77036
rect 1397 77027 1455 77033
rect 1397 77024 1409 77027
rect 1360 76996 1409 77024
rect 1360 76984 1366 76996
rect 1397 76993 1409 76996
rect 1443 76993 1455 77027
rect 1397 76987 1455 76993
rect 1486 76984 1492 77036
rect 1544 77024 1550 77036
rect 2041 77027 2099 77033
rect 2041 77024 2053 77027
rect 1544 76996 2053 77024
rect 1544 76984 1550 76996
rect 2041 76993 2053 76996
rect 2087 76993 2099 77027
rect 2041 76987 2099 76993
rect 2685 77027 2743 77033
rect 2685 76993 2697 77027
rect 2731 77024 2743 77027
rect 3050 77024 3056 77036
rect 2731 76996 3056 77024
rect 2731 76993 2743 76996
rect 2685 76987 2743 76993
rect 3050 76984 3056 76996
rect 3108 76984 3114 77036
rect 8294 76984 8300 77036
rect 8352 77024 8358 77036
rect 9125 77027 9183 77033
rect 9125 77024 9137 77027
rect 8352 76996 9137 77024
rect 8352 76984 8358 76996
rect 9125 76993 9137 76996
rect 9171 76993 9183 77027
rect 9125 76987 9183 76993
rect 9674 76984 9680 77036
rect 9732 77024 9738 77036
rect 9861 77027 9919 77033
rect 9861 77024 9873 77027
rect 9732 76996 9873 77024
rect 9732 76984 9738 76996
rect 9861 76993 9873 76996
rect 9907 76993 9919 77027
rect 9861 76987 9919 76993
rect 1578 76820 1584 76832
rect 1539 76792 1584 76820
rect 1578 76780 1584 76792
rect 1636 76780 1642 76832
rect 2222 76820 2228 76832
rect 2183 76792 2228 76820
rect 2222 76780 2228 76792
rect 2280 76780 2286 76832
rect 2869 76823 2927 76829
rect 2869 76789 2881 76823
rect 2915 76820 2927 76823
rect 3602 76820 3608 76832
rect 2915 76792 3608 76820
rect 2915 76789 2927 76792
rect 2869 76783 2927 76789
rect 3602 76780 3608 76792
rect 3660 76780 3666 76832
rect 10042 76820 10048 76832
rect 10003 76792 10048 76820
rect 10042 76780 10048 76792
rect 10100 76780 10106 76832
rect 1104 76730 10856 76752
rect 1104 76678 2582 76730
rect 2634 76678 2646 76730
rect 2698 76678 2710 76730
rect 2762 76678 2774 76730
rect 2826 76678 2838 76730
rect 2890 76678 5845 76730
rect 5897 76678 5909 76730
rect 5961 76678 5973 76730
rect 6025 76678 6037 76730
rect 6089 76678 6101 76730
rect 6153 76678 9109 76730
rect 9161 76678 9173 76730
rect 9225 76678 9237 76730
rect 9289 76678 9301 76730
rect 9353 76678 9365 76730
rect 9417 76678 10856 76730
rect 1104 76656 10856 76678
rect 10045 76619 10103 76625
rect 10045 76585 10057 76619
rect 10091 76616 10103 76619
rect 10965 76619 11023 76625
rect 10965 76616 10977 76619
rect 10091 76588 10977 76616
rect 10091 76585 10103 76588
rect 10045 76579 10103 76585
rect 10965 76585 10977 76588
rect 11011 76585 11023 76619
rect 10965 76579 11023 76585
rect 1394 76412 1400 76424
rect 1355 76384 1400 76412
rect 1394 76372 1400 76384
rect 1452 76372 1458 76424
rect 9766 76372 9772 76424
rect 9824 76412 9830 76424
rect 9861 76415 9919 76421
rect 9861 76412 9873 76415
rect 9824 76384 9873 76412
rect 9824 76372 9830 76384
rect 9861 76381 9873 76384
rect 9907 76381 9919 76415
rect 9861 76375 9919 76381
rect 1486 76236 1492 76288
rect 1544 76276 1550 76288
rect 1581 76279 1639 76285
rect 1581 76276 1593 76279
rect 1544 76248 1593 76276
rect 1544 76236 1550 76248
rect 1581 76245 1593 76248
rect 1627 76245 1639 76279
rect 1581 76239 1639 76245
rect 1104 76186 10856 76208
rect 1104 76134 4213 76186
rect 4265 76134 4277 76186
rect 4329 76134 4341 76186
rect 4393 76134 4405 76186
rect 4457 76134 4469 76186
rect 4521 76134 7477 76186
rect 7529 76134 7541 76186
rect 7593 76134 7605 76186
rect 7657 76134 7669 76186
rect 7721 76134 7733 76186
rect 7785 76134 10856 76186
rect 1104 76112 10856 76134
rect 1581 76075 1639 76081
rect 1581 76041 1593 76075
rect 1627 76072 1639 76075
rect 3050 76072 3056 76084
rect 1627 76044 3056 76072
rect 1627 76041 1639 76044
rect 1581 76035 1639 76041
rect 3050 76032 3056 76044
rect 3108 76032 3114 76084
rect 1302 75896 1308 75948
rect 1360 75936 1366 75948
rect 1397 75939 1455 75945
rect 1397 75936 1409 75939
rect 1360 75908 1409 75936
rect 1360 75896 1366 75908
rect 1397 75905 1409 75908
rect 1443 75905 1455 75939
rect 1397 75899 1455 75905
rect 9861 75939 9919 75945
rect 9861 75905 9873 75939
rect 9907 75905 9919 75939
rect 9861 75899 9919 75905
rect 6270 75828 6276 75880
rect 6328 75868 6334 75880
rect 9876 75868 9904 75899
rect 6328 75840 9904 75868
rect 6328 75828 6334 75840
rect 10042 75732 10048 75744
rect 10003 75704 10048 75732
rect 10042 75692 10048 75704
rect 10100 75692 10106 75744
rect 1104 75642 10856 75664
rect 1104 75590 2582 75642
rect 2634 75590 2646 75642
rect 2698 75590 2710 75642
rect 2762 75590 2774 75642
rect 2826 75590 2838 75642
rect 2890 75590 5845 75642
rect 5897 75590 5909 75642
rect 5961 75590 5973 75642
rect 6025 75590 6037 75642
rect 6089 75590 6101 75642
rect 6153 75590 9109 75642
rect 9161 75590 9173 75642
rect 9225 75590 9237 75642
rect 9289 75590 9301 75642
rect 9353 75590 9365 75642
rect 9417 75590 10856 75642
rect 1104 75568 10856 75590
rect 1581 75463 1639 75469
rect 1581 75429 1593 75463
rect 1627 75460 1639 75463
rect 3142 75460 3148 75472
rect 1627 75432 3148 75460
rect 1627 75429 1639 75432
rect 1581 75423 1639 75429
rect 3142 75420 3148 75432
rect 3200 75420 3206 75472
rect 1394 75324 1400 75336
rect 1355 75296 1400 75324
rect 1394 75284 1400 75296
rect 1452 75284 1458 75336
rect 2038 75324 2044 75336
rect 1999 75296 2044 75324
rect 2038 75284 2044 75296
rect 2096 75284 2102 75336
rect 9858 75324 9864 75336
rect 9819 75296 9864 75324
rect 9858 75284 9864 75296
rect 9916 75284 9922 75336
rect 2225 75191 2283 75197
rect 2225 75157 2237 75191
rect 2271 75188 2283 75191
rect 2958 75188 2964 75200
rect 2271 75160 2964 75188
rect 2271 75157 2283 75160
rect 2225 75151 2283 75157
rect 2958 75148 2964 75160
rect 3016 75148 3022 75200
rect 10042 75188 10048 75200
rect 10003 75160 10048 75188
rect 10042 75148 10048 75160
rect 10100 75148 10106 75200
rect 1104 75098 10856 75120
rect 1104 75046 4213 75098
rect 4265 75046 4277 75098
rect 4329 75046 4341 75098
rect 4393 75046 4405 75098
rect 4457 75046 4469 75098
rect 4521 75046 7477 75098
rect 7529 75046 7541 75098
rect 7593 75046 7605 75098
rect 7657 75046 7669 75098
rect 7721 75046 7733 75098
rect 7785 75046 10856 75098
rect 1104 75024 10856 75046
rect 2961 74987 3019 74993
rect 1596 74956 2912 74984
rect 1596 74925 1624 74956
rect 1581 74919 1639 74925
rect 1581 74885 1593 74919
rect 1627 74885 1639 74919
rect 1581 74879 1639 74885
rect 1670 74876 1676 74928
rect 1728 74916 1734 74928
rect 1728 74888 1773 74916
rect 1728 74876 1734 74888
rect 2222 74876 2228 74928
rect 2280 74916 2286 74928
rect 2685 74919 2743 74925
rect 2685 74916 2697 74919
rect 2280 74888 2697 74916
rect 2280 74876 2286 74888
rect 2685 74885 2697 74888
rect 2731 74885 2743 74919
rect 2884 74916 2912 74956
rect 2961 74953 2973 74987
rect 3007 74984 3019 74987
rect 5534 74984 5540 74996
rect 3007 74956 5540 74984
rect 3007 74953 3019 74956
rect 2961 74947 3019 74953
rect 5534 74944 5540 74956
rect 5592 74944 5598 74996
rect 6546 74916 6552 74928
rect 2884 74888 6552 74916
rect 2685 74879 2743 74885
rect 6546 74876 6552 74888
rect 6604 74876 6610 74928
rect 1397 74851 1455 74857
rect 1397 74817 1409 74851
rect 1443 74848 1455 74851
rect 1765 74851 1823 74857
rect 1443 74820 1716 74848
rect 1443 74817 1455 74820
rect 1397 74811 1455 74817
rect 1688 74792 1716 74820
rect 1765 74817 1777 74851
rect 1811 74848 1823 74851
rect 2130 74848 2136 74860
rect 1811 74820 2136 74848
rect 1811 74817 1823 74820
rect 1765 74811 1823 74817
rect 2130 74808 2136 74820
rect 2188 74808 2194 74860
rect 2409 74851 2467 74857
rect 2409 74817 2421 74851
rect 2455 74817 2467 74851
rect 2590 74848 2596 74860
rect 2551 74820 2596 74848
rect 2409 74811 2467 74817
rect 1670 74740 1676 74792
rect 1728 74740 1734 74792
rect 2424 74780 2452 74811
rect 2590 74808 2596 74820
rect 2648 74808 2654 74860
rect 2777 74851 2835 74857
rect 2777 74817 2789 74851
rect 2823 74848 2835 74851
rect 3694 74848 3700 74860
rect 2823 74820 3700 74848
rect 2823 74817 2835 74820
rect 2777 74811 2835 74817
rect 3694 74808 3700 74820
rect 3752 74808 3758 74860
rect 3510 74780 3516 74792
rect 2424 74752 3516 74780
rect 3510 74740 3516 74752
rect 3568 74740 3574 74792
rect 1118 74672 1124 74724
rect 1176 74712 1182 74724
rect 2590 74712 2596 74724
rect 1176 74684 2596 74712
rect 1176 74672 1182 74684
rect 2590 74672 2596 74684
rect 2648 74672 2654 74724
rect 1949 74647 2007 74653
rect 1949 74613 1961 74647
rect 1995 74644 2007 74647
rect 6270 74644 6276 74656
rect 1995 74616 6276 74644
rect 1995 74613 2007 74616
rect 1949 74607 2007 74613
rect 6270 74604 6276 74616
rect 6328 74604 6334 74656
rect 1104 74554 10856 74576
rect 1104 74502 2582 74554
rect 2634 74502 2646 74554
rect 2698 74502 2710 74554
rect 2762 74502 2774 74554
rect 2826 74502 2838 74554
rect 2890 74502 5845 74554
rect 5897 74502 5909 74554
rect 5961 74502 5973 74554
rect 6025 74502 6037 74554
rect 6089 74502 6101 74554
rect 6153 74502 9109 74554
rect 9161 74502 9173 74554
rect 9225 74502 9237 74554
rect 9289 74502 9301 74554
rect 9353 74502 9365 74554
rect 9417 74502 10856 74554
rect 1104 74480 10856 74502
rect 1949 74443 2007 74449
rect 1949 74409 1961 74443
rect 1995 74440 2007 74443
rect 9858 74440 9864 74452
rect 1995 74412 9864 74440
rect 1995 74409 2007 74412
rect 1949 74403 2007 74409
rect 9858 74400 9864 74412
rect 9916 74400 9922 74452
rect 2961 74375 3019 74381
rect 2961 74341 2973 74375
rect 3007 74372 3019 74375
rect 9674 74372 9680 74384
rect 3007 74344 9680 74372
rect 3007 74341 3019 74344
rect 2961 74335 3019 74341
rect 9674 74332 9680 74344
rect 9732 74332 9738 74384
rect 1578 74264 1584 74316
rect 1636 74304 1642 74316
rect 5626 74304 5632 74316
rect 1636 74276 1716 74304
rect 1636 74264 1642 74276
rect 1688 74245 1716 74276
rect 3436 74276 5632 74304
rect 1397 74239 1455 74245
rect 1397 74205 1409 74239
rect 1443 74205 1455 74239
rect 1397 74199 1455 74205
rect 1673 74239 1731 74245
rect 1673 74205 1685 74239
rect 1719 74205 1731 74239
rect 1673 74199 1731 74205
rect 1765 74239 1823 74245
rect 1765 74205 1777 74239
rect 1811 74236 1823 74239
rect 2130 74236 2136 74248
rect 1811 74208 2136 74236
rect 1811 74205 1823 74208
rect 1765 74199 1823 74205
rect 1412 74100 1440 74199
rect 2130 74196 2136 74208
rect 2188 74196 2194 74248
rect 2409 74239 2467 74245
rect 2409 74205 2421 74239
rect 2455 74205 2467 74239
rect 2682 74236 2688 74248
rect 2643 74208 2688 74236
rect 2409 74199 2467 74205
rect 1578 74168 1584 74180
rect 1539 74140 1584 74168
rect 1578 74128 1584 74140
rect 1636 74128 1642 74180
rect 2424 74168 2452 74199
rect 2682 74196 2688 74208
rect 2740 74196 2746 74248
rect 2774 74196 2780 74248
rect 2832 74236 2838 74248
rect 2832 74208 2877 74236
rect 2832 74196 2838 74208
rect 1688 74140 2452 74168
rect 2593 74171 2651 74177
rect 1688 74112 1716 74140
rect 2593 74137 2605 74171
rect 2639 74168 2651 74171
rect 3326 74168 3332 74180
rect 2639 74140 3332 74168
rect 2639 74137 2651 74140
rect 2593 74131 2651 74137
rect 3326 74128 3332 74140
rect 3384 74128 3390 74180
rect 1670 74100 1676 74112
rect 1412 74072 1676 74100
rect 1670 74060 1676 74072
rect 1728 74060 1734 74112
rect 2498 74060 2504 74112
rect 2556 74100 2562 74112
rect 3436 74100 3464 74276
rect 5626 74264 5632 74276
rect 5684 74264 5690 74316
rect 3786 74236 3792 74248
rect 3747 74208 3792 74236
rect 3786 74196 3792 74208
rect 3844 74196 3850 74248
rect 3970 74196 3976 74248
rect 4028 74236 4034 74248
rect 4798 74236 4804 74248
rect 4028 74208 4804 74236
rect 4028 74196 4034 74208
rect 4798 74196 4804 74208
rect 4856 74196 4862 74248
rect 9858 74236 9864 74248
rect 9819 74208 9864 74236
rect 9858 74196 9864 74208
rect 9916 74196 9922 74248
rect 3694 74128 3700 74180
rect 3752 74168 3758 74180
rect 4982 74168 4988 74180
rect 3752 74140 4988 74168
rect 3752 74128 3758 74140
rect 4982 74128 4988 74140
rect 5040 74128 5046 74180
rect 2556 74072 3464 74100
rect 3973 74103 4031 74109
rect 2556 74060 2562 74072
rect 3973 74069 3985 74103
rect 4019 74100 4031 74103
rect 4062 74100 4068 74112
rect 4019 74072 4068 74100
rect 4019 74069 4031 74072
rect 3973 74063 4031 74069
rect 4062 74060 4068 74072
rect 4120 74060 4126 74112
rect 10042 74100 10048 74112
rect 10003 74072 10048 74100
rect 10042 74060 10048 74072
rect 10100 74060 10106 74112
rect 1104 74010 10856 74032
rect 1104 73958 4213 74010
rect 4265 73958 4277 74010
rect 4329 73958 4341 74010
rect 4393 73958 4405 74010
rect 4457 73958 4469 74010
rect 4521 73958 7477 74010
rect 7529 73958 7541 74010
rect 7593 73958 7605 74010
rect 7657 73958 7669 74010
rect 7721 73958 7733 74010
rect 7785 73958 10856 74010
rect 1104 73936 10856 73958
rect 2498 73856 2504 73908
rect 2556 73896 2562 73908
rect 3053 73899 3111 73905
rect 2556 73868 2728 73896
rect 2556 73856 2562 73868
rect 1486 73788 1492 73840
rect 1544 73828 1550 73840
rect 2700 73837 2728 73868
rect 3053 73865 3065 73899
rect 3099 73896 3111 73899
rect 4065 73899 4123 73905
rect 3099 73868 4016 73896
rect 3099 73865 3111 73868
rect 3053 73859 3111 73865
rect 1673 73831 1731 73837
rect 1673 73828 1685 73831
rect 1544 73800 1685 73828
rect 1544 73788 1550 73800
rect 1673 73797 1685 73800
rect 1719 73797 1731 73831
rect 1673 73791 1731 73797
rect 2685 73831 2743 73837
rect 2685 73797 2697 73831
rect 2731 73797 2743 73831
rect 2685 73791 2743 73797
rect 2777 73831 2835 73837
rect 2777 73797 2789 73831
rect 2823 73828 2835 73831
rect 2958 73828 2964 73840
rect 2823 73800 2964 73828
rect 2823 73797 2835 73800
rect 2777 73791 2835 73797
rect 2958 73788 2964 73800
rect 3016 73788 3022 73840
rect 3602 73788 3608 73840
rect 3660 73828 3666 73840
rect 3789 73831 3847 73837
rect 3789 73828 3801 73831
rect 3660 73800 3801 73828
rect 3660 73788 3666 73800
rect 3789 73797 3801 73800
rect 3835 73797 3847 73831
rect 3789 73791 3847 73797
rect 1397 73763 1455 73769
rect 1397 73729 1409 73763
rect 1443 73760 1455 73763
rect 1581 73763 1639 73769
rect 1443 73732 1532 73760
rect 1443 73729 1455 73732
rect 1397 73723 1455 73729
rect 1504 73636 1532 73732
rect 1581 73729 1593 73763
rect 1627 73729 1639 73763
rect 1581 73723 1639 73729
rect 1765 73763 1823 73769
rect 1765 73729 1777 73763
rect 1811 73760 1823 73763
rect 2130 73760 2136 73772
rect 1811 73732 2136 73760
rect 1811 73729 1823 73732
rect 1765 73723 1823 73729
rect 1596 73692 1624 73723
rect 2130 73720 2136 73732
rect 2188 73720 2194 73772
rect 2406 73720 2412 73772
rect 2464 73760 2470 73772
rect 2501 73763 2559 73769
rect 2501 73760 2513 73763
rect 2464 73732 2513 73760
rect 2464 73720 2470 73732
rect 2501 73729 2513 73732
rect 2547 73729 2559 73763
rect 2501 73723 2559 73729
rect 2869 73763 2927 73769
rect 2869 73729 2881 73763
rect 2915 73760 2927 73763
rect 3510 73760 3516 73772
rect 2915 73732 3004 73760
rect 3471 73732 3516 73760
rect 2915 73729 2927 73732
rect 2869 73723 2927 73729
rect 2148 73692 2176 73720
rect 2976 73704 3004 73732
rect 3510 73720 3516 73732
rect 3568 73720 3574 73772
rect 3697 73763 3755 73769
rect 3697 73729 3709 73763
rect 3743 73729 3755 73763
rect 3697 73723 3755 73729
rect 3881 73763 3939 73769
rect 3881 73729 3893 73763
rect 3927 73729 3939 73763
rect 3881 73723 3939 73729
rect 2774 73692 2780 73704
rect 1596 73664 1808 73692
rect 2148 73664 2780 73692
rect 1486 73584 1492 73636
rect 1544 73624 1550 73636
rect 1670 73624 1676 73636
rect 1544 73596 1676 73624
rect 1544 73584 1550 73596
rect 1670 73584 1676 73596
rect 1728 73584 1734 73636
rect 474 73516 480 73568
rect 532 73556 538 73568
rect 1780 73556 1808 73664
rect 2774 73652 2780 73664
rect 2832 73652 2838 73704
rect 2958 73652 2964 73704
rect 3016 73652 3022 73704
rect 3712 73624 3740 73723
rect 3786 73652 3792 73704
rect 3844 73692 3850 73704
rect 3896 73692 3924 73723
rect 3844 73664 3924 73692
rect 3988 73692 4016 73868
rect 4065 73865 4077 73899
rect 4111 73896 4123 73899
rect 5077 73899 5135 73905
rect 4111 73868 5028 73896
rect 4111 73865 4123 73868
rect 4065 73859 4123 73865
rect 4706 73788 4712 73840
rect 4764 73828 4770 73840
rect 5000 73828 5028 73868
rect 5077 73865 5089 73899
rect 5123 73896 5135 73899
rect 8294 73896 8300 73908
rect 5123 73868 8300 73896
rect 5123 73865 5135 73868
rect 5077 73859 5135 73865
rect 8294 73856 8300 73868
rect 8352 73856 8358 73908
rect 9766 73828 9772 73840
rect 4764 73800 4809 73828
rect 5000 73800 9772 73828
rect 4764 73788 4770 73800
rect 9766 73788 9772 73800
rect 9824 73788 9830 73840
rect 4522 73720 4528 73772
rect 4580 73769 4586 73772
rect 4798 73769 4804 73772
rect 4580 73763 4603 73769
rect 4591 73729 4603 73763
rect 4580 73723 4603 73729
rect 4797 73723 4804 73769
rect 4856 73760 4862 73772
rect 4982 73769 4988 73772
rect 4939 73763 4988 73769
rect 4856 73732 4897 73760
rect 4580 73720 4586 73723
rect 4798 73720 4804 73723
rect 4856 73720 4862 73732
rect 4939 73729 4951 73763
rect 4985 73729 4988 73763
rect 4939 73723 4988 73729
rect 4982 73720 4988 73723
rect 5040 73720 5046 73772
rect 9861 73763 9919 73769
rect 9861 73729 9873 73763
rect 9907 73729 9919 73763
rect 9861 73723 9919 73729
rect 9876 73692 9904 73723
rect 3988 73664 9904 73692
rect 3844 73652 3850 73664
rect 4982 73624 4988 73636
rect 3712 73596 4988 73624
rect 4982 73584 4988 73596
rect 5040 73584 5046 73636
rect 532 73528 1808 73556
rect 1949 73559 2007 73565
rect 532 73516 538 73528
rect 1949 73525 1961 73559
rect 1995 73556 2007 73559
rect 9858 73556 9864 73568
rect 1995 73528 9864 73556
rect 1995 73525 2007 73528
rect 1949 73519 2007 73525
rect 9858 73516 9864 73528
rect 9916 73516 9922 73568
rect 10042 73556 10048 73568
rect 10003 73528 10048 73556
rect 10042 73516 10048 73528
rect 10100 73516 10106 73568
rect 1104 73466 10856 73488
rect 1104 73414 2582 73466
rect 2634 73414 2646 73466
rect 2698 73414 2710 73466
rect 2762 73414 2774 73466
rect 2826 73414 2838 73466
rect 2890 73414 5845 73466
rect 5897 73414 5909 73466
rect 5961 73414 5973 73466
rect 6025 73414 6037 73466
rect 6089 73414 6101 73466
rect 6153 73414 9109 73466
rect 9161 73414 9173 73466
rect 9225 73414 9237 73466
rect 9289 73414 9301 73466
rect 9353 73414 9365 73466
rect 9417 73414 10856 73466
rect 1104 73392 10856 73414
rect 1578 73312 1584 73364
rect 1636 73352 1642 73364
rect 4798 73352 4804 73364
rect 1636 73324 4804 73352
rect 1636 73312 1642 73324
rect 4798 73312 4804 73324
rect 4856 73312 4862 73364
rect 3053 73287 3111 73293
rect 3053 73253 3065 73287
rect 3099 73253 3111 73287
rect 3053 73247 3111 73253
rect 1397 73151 1455 73157
rect 1397 73117 1409 73151
rect 1443 73148 1455 73151
rect 1486 73148 1492 73160
rect 1443 73120 1492 73148
rect 1443 73117 1455 73120
rect 1397 73111 1455 73117
rect 1486 73108 1492 73120
rect 1544 73108 1550 73160
rect 1670 73148 1676 73160
rect 1631 73120 1676 73148
rect 1670 73108 1676 73120
rect 1728 73108 1734 73160
rect 1765 73151 1823 73157
rect 1765 73117 1777 73151
rect 1811 73148 1823 73151
rect 2130 73148 2136 73160
rect 1811 73120 2136 73148
rect 1811 73117 1823 73120
rect 1765 73111 1823 73117
rect 2130 73108 2136 73120
rect 2188 73108 2194 73160
rect 2406 73108 2412 73160
rect 2464 73148 2470 73160
rect 2501 73151 2559 73157
rect 2501 73148 2513 73151
rect 2464 73120 2513 73148
rect 2464 73108 2470 73120
rect 2501 73117 2513 73120
rect 2547 73117 2559 73151
rect 2866 73148 2872 73160
rect 2827 73120 2872 73148
rect 2501 73111 2559 73117
rect 2866 73108 2872 73120
rect 2924 73108 2930 73160
rect 2958 73108 2964 73160
rect 3016 73108 3022 73160
rect 3068 73148 3096 73247
rect 3510 73176 3516 73228
rect 3568 73216 3574 73228
rect 4522 73216 4528 73228
rect 3568 73188 4528 73216
rect 3568 73176 3574 73188
rect 4522 73176 4528 73188
rect 4580 73176 4586 73228
rect 9861 73151 9919 73157
rect 9861 73148 9873 73151
rect 3068 73120 9873 73148
rect 9861 73117 9873 73120
rect 9907 73117 9919 73151
rect 9861 73111 9919 73117
rect 1578 73080 1584 73092
rect 1539 73052 1584 73080
rect 1578 73040 1584 73052
rect 1636 73040 1642 73092
rect 2685 73083 2743 73089
rect 2685 73080 2697 73083
rect 1872 73052 2697 73080
rect 842 72972 848 73024
rect 900 73012 906 73024
rect 1872 73012 1900 73052
rect 2685 73049 2697 73052
rect 2731 73049 2743 73083
rect 2685 73043 2743 73049
rect 2777 73083 2835 73089
rect 2777 73049 2789 73083
rect 2823 73080 2835 73083
rect 2976 73080 3004 73108
rect 11057 73083 11115 73089
rect 11057 73080 11069 73083
rect 2823 73052 3004 73080
rect 3160 73052 11069 73080
rect 2823 73049 2835 73052
rect 2777 73043 2835 73049
rect 900 72984 1900 73012
rect 1949 73015 2007 73021
rect 900 72972 906 72984
rect 1949 72981 1961 73015
rect 1995 73012 2007 73015
rect 3160 73012 3188 73052
rect 11057 73049 11069 73052
rect 11103 73049 11115 73083
rect 11057 73043 11115 73049
rect 10042 73012 10048 73024
rect 1995 72984 3188 73012
rect 10003 72984 10048 73012
rect 1995 72981 2007 72984
rect 1949 72975 2007 72981
rect 10042 72972 10048 72984
rect 10100 72972 10106 73024
rect 1104 72922 10856 72944
rect 1104 72870 4213 72922
rect 4265 72870 4277 72922
rect 4329 72870 4341 72922
rect 4393 72870 4405 72922
rect 4457 72870 4469 72922
rect 4521 72870 7477 72922
rect 7529 72870 7541 72922
rect 7593 72870 7605 72922
rect 7657 72870 7669 72922
rect 7721 72870 7733 72922
rect 7785 72870 10856 72922
rect 1104 72848 10856 72870
rect 1486 72700 1492 72752
rect 1544 72740 1550 72752
rect 1544 72712 4292 72740
rect 1544 72700 1550 72712
rect 1394 72672 1400 72684
rect 1355 72644 1400 72672
rect 1394 72632 1400 72644
rect 1452 72632 1458 72684
rect 2038 72672 2044 72684
rect 1999 72644 2044 72672
rect 2038 72632 2044 72644
rect 2096 72632 2102 72684
rect 2130 72632 2136 72684
rect 2188 72672 2194 72684
rect 4264 72681 4292 72712
rect 2961 72675 3019 72681
rect 2961 72672 2973 72675
rect 2188 72644 2973 72672
rect 2188 72632 2194 72644
rect 2961 72641 2973 72644
rect 3007 72641 3019 72675
rect 2961 72635 3019 72641
rect 4249 72675 4307 72681
rect 4249 72641 4261 72675
rect 4295 72641 4307 72675
rect 4249 72635 4307 72641
rect 1578 72564 1584 72616
rect 1636 72564 1642 72616
rect 2685 72607 2743 72613
rect 2685 72573 2697 72607
rect 2731 72604 2743 72607
rect 3786 72604 3792 72616
rect 2731 72576 3792 72604
rect 2731 72573 2743 72576
rect 2685 72567 2743 72573
rect 3786 72564 3792 72576
rect 3844 72564 3850 72616
rect 3970 72604 3976 72616
rect 3931 72576 3976 72604
rect 3970 72564 3976 72576
rect 4028 72564 4034 72616
rect 1596 72536 1624 72564
rect 7006 72536 7012 72548
rect 1596 72508 7012 72536
rect 7006 72496 7012 72508
rect 7064 72496 7070 72548
rect 1581 72471 1639 72477
rect 1581 72437 1593 72471
rect 1627 72468 1639 72471
rect 1670 72468 1676 72480
rect 1627 72440 1676 72468
rect 1627 72437 1639 72440
rect 1581 72431 1639 72437
rect 1670 72428 1676 72440
rect 1728 72428 1734 72480
rect 2225 72471 2283 72477
rect 2225 72437 2237 72471
rect 2271 72468 2283 72471
rect 2314 72468 2320 72480
rect 2271 72440 2320 72468
rect 2271 72437 2283 72440
rect 2225 72431 2283 72437
rect 2314 72428 2320 72440
rect 2372 72428 2378 72480
rect 2498 72428 2504 72480
rect 2556 72468 2562 72480
rect 5718 72468 5724 72480
rect 2556 72440 5724 72468
rect 2556 72428 2562 72440
rect 5718 72428 5724 72440
rect 5776 72428 5782 72480
rect 1104 72378 10856 72400
rect 1104 72326 2582 72378
rect 2634 72326 2646 72378
rect 2698 72326 2710 72378
rect 2762 72326 2774 72378
rect 2826 72326 2838 72378
rect 2890 72326 5845 72378
rect 5897 72326 5909 72378
rect 5961 72326 5973 72378
rect 6025 72326 6037 72378
rect 6089 72326 6101 72378
rect 6153 72326 9109 72378
rect 9161 72326 9173 72378
rect 9225 72326 9237 72378
rect 9289 72326 9301 72378
rect 9353 72326 9365 72378
rect 9417 72326 10856 72378
rect 1104 72304 10856 72326
rect 1581 72267 1639 72273
rect 1581 72233 1593 72267
rect 1627 72264 1639 72267
rect 3602 72264 3608 72276
rect 1627 72236 3608 72264
rect 1627 72233 1639 72236
rect 1581 72227 1639 72233
rect 3602 72224 3608 72236
rect 3660 72224 3666 72276
rect 2498 72156 2504 72208
rect 2556 72156 2562 72208
rect 4341 72199 4399 72205
rect 4341 72165 4353 72199
rect 4387 72165 4399 72199
rect 4341 72159 4399 72165
rect 2516 72128 2544 72156
rect 3142 72128 3148 72140
rect 2516 72100 2728 72128
rect 1394 72060 1400 72072
rect 1355 72032 1400 72060
rect 1394 72020 1400 72032
rect 1452 72020 1458 72072
rect 2406 72020 2412 72072
rect 2464 72060 2470 72072
rect 2700 72069 2728 72100
rect 2792 72100 3148 72128
rect 2792 72069 2820 72100
rect 3142 72088 3148 72100
rect 3200 72088 3206 72140
rect 3712 72100 4200 72128
rect 2501 72063 2559 72069
rect 2501 72060 2513 72063
rect 2464 72032 2513 72060
rect 2464 72020 2470 72032
rect 2501 72029 2513 72032
rect 2547 72029 2559 72063
rect 2501 72023 2559 72029
rect 2685 72063 2743 72069
rect 2685 72029 2697 72063
rect 2731 72029 2743 72063
rect 2685 72023 2743 72029
rect 2777 72063 2835 72069
rect 2777 72029 2789 72063
rect 2823 72029 2835 72063
rect 2777 72023 2835 72029
rect 2869 72063 2927 72069
rect 2869 72029 2881 72063
rect 2915 72060 2927 72063
rect 2958 72060 2964 72072
rect 2915 72032 2964 72060
rect 2915 72029 2927 72032
rect 2869 72023 2927 72029
rect 2516 71924 2544 72023
rect 2958 72020 2964 72032
rect 3016 72060 3022 72072
rect 3712 72060 3740 72100
rect 3016 72032 3740 72060
rect 3789 72063 3847 72069
rect 3016 72020 3022 72032
rect 3789 72029 3801 72063
rect 3835 72060 3847 72063
rect 3878 72060 3884 72072
rect 3835 72032 3884 72060
rect 3835 72029 3847 72032
rect 3789 72023 3847 72029
rect 3804 71992 3832 72023
rect 3878 72020 3884 72032
rect 3936 72020 3942 72072
rect 4062 72060 4068 72072
rect 4023 72032 4068 72060
rect 4062 72020 4068 72032
rect 4120 72020 4126 72072
rect 4172 72069 4200 72100
rect 4157 72063 4215 72069
rect 4157 72029 4169 72063
rect 4203 72029 4215 72063
rect 4356 72060 4384 72159
rect 9861 72063 9919 72069
rect 9861 72060 9873 72063
rect 4356 72032 9873 72060
rect 4157 72023 4215 72029
rect 9861 72029 9873 72032
rect 9907 72029 9919 72063
rect 9861 72023 9919 72029
rect 2884 71964 3832 71992
rect 3973 71995 4031 72001
rect 2884 71936 2912 71964
rect 3973 71961 3985 71995
rect 4019 71992 4031 71995
rect 6454 71992 6460 72004
rect 4019 71964 6460 71992
rect 4019 71961 4031 71964
rect 3973 71955 4031 71961
rect 6454 71952 6460 71964
rect 6512 71952 6518 72004
rect 2866 71924 2872 71936
rect 2516 71896 2872 71924
rect 2866 71884 2872 71896
rect 2924 71884 2930 71936
rect 3053 71927 3111 71933
rect 3053 71893 3065 71927
rect 3099 71924 3111 71927
rect 9858 71924 9864 71936
rect 3099 71896 9864 71924
rect 3099 71893 3111 71896
rect 3053 71887 3111 71893
rect 9858 71884 9864 71896
rect 9916 71884 9922 71936
rect 10042 71924 10048 71936
rect 10003 71896 10048 71924
rect 10042 71884 10048 71896
rect 10100 71884 10106 71936
rect 1104 71834 10856 71856
rect 1104 71782 4213 71834
rect 4265 71782 4277 71834
rect 4329 71782 4341 71834
rect 4393 71782 4405 71834
rect 4457 71782 4469 71834
rect 4521 71782 7477 71834
rect 7529 71782 7541 71834
rect 7593 71782 7605 71834
rect 7657 71782 7669 71834
rect 7721 71782 7733 71834
rect 7785 71782 10856 71834
rect 1104 71760 10856 71782
rect 4614 71720 4620 71732
rect 2148 71692 4620 71720
rect 1394 71584 1400 71596
rect 1355 71556 1400 71584
rect 1394 71544 1400 71556
rect 1452 71544 1458 71596
rect 2041 71587 2099 71593
rect 2041 71553 2053 71587
rect 2087 71553 2099 71587
rect 2148 71584 2176 71692
rect 4614 71680 4620 71692
rect 4672 71680 4678 71732
rect 2314 71652 2320 71664
rect 2275 71624 2320 71652
rect 2314 71612 2320 71624
rect 2372 71612 2378 71664
rect 2225 71587 2283 71593
rect 2225 71584 2237 71587
rect 2148 71556 2237 71584
rect 2041 71547 2099 71553
rect 2225 71553 2237 71556
rect 2271 71553 2283 71587
rect 2225 71547 2283 71553
rect 2409 71587 2467 71593
rect 2409 71553 2421 71587
rect 2455 71584 2467 71587
rect 2958 71584 2964 71596
rect 2455 71556 2964 71584
rect 2455 71553 2467 71556
rect 2409 71547 2467 71553
rect 2056 71516 2084 71547
rect 2958 71544 2964 71556
rect 3016 71584 3022 71596
rect 3605 71587 3663 71593
rect 3605 71584 3617 71587
rect 3016 71556 3617 71584
rect 3016 71544 3022 71556
rect 3605 71553 3617 71556
rect 3651 71553 3663 71587
rect 3605 71547 3663 71553
rect 3786 71544 3792 71596
rect 3844 71584 3850 71596
rect 3881 71587 3939 71593
rect 3881 71584 3893 71587
rect 3844 71556 3893 71584
rect 3844 71544 3850 71556
rect 3881 71553 3893 71556
rect 3927 71553 3939 71587
rect 9858 71584 9864 71596
rect 9819 71556 9864 71584
rect 3881 71547 3939 71553
rect 9858 71544 9864 71556
rect 9916 71544 9922 71596
rect 2866 71516 2872 71528
rect 2056 71488 2872 71516
rect 2866 71476 2872 71488
rect 2924 71476 2930 71528
rect 1581 71383 1639 71389
rect 1581 71349 1593 71383
rect 1627 71380 1639 71383
rect 2498 71380 2504 71392
rect 1627 71352 2504 71380
rect 1627 71349 1639 71352
rect 1581 71343 1639 71349
rect 2498 71340 2504 71352
rect 2556 71340 2562 71392
rect 2593 71383 2651 71389
rect 2593 71349 2605 71383
rect 2639 71380 2651 71383
rect 9858 71380 9864 71392
rect 2639 71352 9864 71380
rect 2639 71349 2651 71352
rect 2593 71343 2651 71349
rect 9858 71340 9864 71352
rect 9916 71340 9922 71392
rect 10042 71380 10048 71392
rect 10003 71352 10048 71380
rect 10042 71340 10048 71352
rect 10100 71340 10106 71392
rect 1104 71290 10856 71312
rect 1104 71238 2582 71290
rect 2634 71238 2646 71290
rect 2698 71238 2710 71290
rect 2762 71238 2774 71290
rect 2826 71238 2838 71290
rect 2890 71238 5845 71290
rect 5897 71238 5909 71290
rect 5961 71238 5973 71290
rect 6025 71238 6037 71290
rect 6089 71238 6101 71290
rect 6153 71238 9109 71290
rect 9161 71238 9173 71290
rect 9225 71238 9237 71290
rect 9289 71238 9301 71290
rect 9353 71238 9365 71290
rect 9417 71238 10856 71290
rect 1104 71216 10856 71238
rect 3789 71043 3847 71049
rect 3789 71009 3801 71043
rect 3835 71040 3847 71043
rect 3970 71040 3976 71052
rect 3835 71012 3976 71040
rect 3835 71009 3847 71012
rect 3789 71003 3847 71009
rect 3970 71000 3976 71012
rect 4028 71000 4034 71052
rect 1394 70972 1400 70984
rect 1355 70944 1400 70972
rect 1394 70932 1400 70944
rect 1452 70932 1458 70984
rect 3878 70932 3884 70984
rect 3936 70972 3942 70984
rect 4065 70975 4123 70981
rect 4065 70972 4077 70975
rect 3936 70944 4077 70972
rect 3936 70932 3942 70944
rect 4065 70941 4077 70944
rect 4111 70941 4123 70975
rect 4065 70935 4123 70941
rect 1581 70839 1639 70845
rect 1581 70805 1593 70839
rect 1627 70836 1639 70839
rect 2406 70836 2412 70848
rect 1627 70808 2412 70836
rect 1627 70805 1639 70808
rect 1581 70799 1639 70805
rect 2406 70796 2412 70808
rect 2464 70796 2470 70848
rect 3694 70796 3700 70848
rect 3752 70836 3758 70848
rect 3878 70836 3884 70848
rect 3752 70808 3884 70836
rect 3752 70796 3758 70808
rect 3878 70796 3884 70808
rect 3936 70796 3942 70848
rect 1104 70746 10856 70768
rect 1104 70694 4213 70746
rect 4265 70694 4277 70746
rect 4329 70694 4341 70746
rect 4393 70694 4405 70746
rect 4457 70694 4469 70746
rect 4521 70694 7477 70746
rect 7529 70694 7541 70746
rect 7593 70694 7605 70746
rect 7657 70694 7669 70746
rect 7721 70694 7733 70746
rect 7785 70694 10856 70746
rect 1104 70672 10856 70694
rect 1581 70635 1639 70641
rect 1581 70601 1593 70635
rect 1627 70632 1639 70635
rect 2038 70632 2044 70644
rect 1627 70604 2044 70632
rect 1627 70601 1639 70604
rect 1581 70595 1639 70601
rect 2038 70592 2044 70604
rect 2096 70592 2102 70644
rect 10045 70635 10103 70641
rect 10045 70601 10057 70635
rect 10091 70632 10103 70635
rect 10686 70632 10692 70644
rect 10091 70604 10692 70632
rect 10091 70601 10103 70604
rect 10045 70595 10103 70601
rect 10686 70592 10692 70604
rect 10744 70592 10750 70644
rect 1394 70496 1400 70508
rect 1355 70468 1400 70496
rect 1394 70456 1400 70468
rect 1452 70456 1458 70508
rect 9858 70496 9864 70508
rect 9819 70468 9864 70496
rect 9858 70456 9864 70468
rect 9916 70456 9922 70508
rect 1104 70202 10856 70224
rect 1104 70150 2582 70202
rect 2634 70150 2646 70202
rect 2698 70150 2710 70202
rect 2762 70150 2774 70202
rect 2826 70150 2838 70202
rect 2890 70150 5845 70202
rect 5897 70150 5909 70202
rect 5961 70150 5973 70202
rect 6025 70150 6037 70202
rect 6089 70150 6101 70202
rect 6153 70150 9109 70202
rect 9161 70150 9173 70202
rect 9225 70150 9237 70202
rect 9289 70150 9301 70202
rect 9353 70150 9365 70202
rect 9417 70150 10856 70202
rect 1104 70128 10856 70150
rect 1394 69884 1400 69896
rect 1355 69856 1400 69884
rect 1394 69844 1400 69856
rect 1452 69844 1458 69896
rect 9861 69887 9919 69893
rect 9861 69853 9873 69887
rect 9907 69884 9919 69887
rect 11057 69887 11115 69893
rect 11057 69884 11069 69887
rect 9907 69856 11069 69884
rect 9907 69853 9919 69856
rect 9861 69847 9919 69853
rect 11057 69853 11069 69856
rect 11103 69853 11115 69887
rect 11057 69847 11115 69853
rect 1581 69751 1639 69757
rect 1581 69717 1593 69751
rect 1627 69748 1639 69751
rect 2314 69748 2320 69760
rect 1627 69720 2320 69748
rect 1627 69717 1639 69720
rect 1581 69711 1639 69717
rect 2314 69708 2320 69720
rect 2372 69708 2378 69760
rect 10042 69748 10048 69760
rect 10003 69720 10048 69748
rect 10042 69708 10048 69720
rect 10100 69708 10106 69760
rect 1104 69658 10856 69680
rect 1104 69606 4213 69658
rect 4265 69606 4277 69658
rect 4329 69606 4341 69658
rect 4393 69606 4405 69658
rect 4457 69606 4469 69658
rect 4521 69606 7477 69658
rect 7529 69606 7541 69658
rect 7593 69606 7605 69658
rect 7657 69606 7669 69658
rect 7721 69606 7733 69658
rect 7785 69606 10856 69658
rect 1104 69584 10856 69606
rect 1394 69408 1400 69420
rect 1355 69380 1400 69408
rect 1394 69368 1400 69380
rect 1452 69368 1458 69420
rect 9861 69411 9919 69417
rect 9861 69377 9873 69411
rect 9907 69408 9919 69411
rect 10965 69411 11023 69417
rect 10965 69408 10977 69411
rect 9907 69380 10977 69408
rect 9907 69377 9919 69380
rect 9861 69371 9919 69377
rect 10965 69377 10977 69380
rect 11011 69377 11023 69411
rect 10965 69371 11023 69377
rect 1581 69207 1639 69213
rect 1581 69173 1593 69207
rect 1627 69204 1639 69207
rect 1762 69204 1768 69216
rect 1627 69176 1768 69204
rect 1627 69173 1639 69176
rect 1581 69167 1639 69173
rect 1762 69164 1768 69176
rect 1820 69164 1826 69216
rect 10042 69204 10048 69216
rect 10003 69176 10048 69204
rect 10042 69164 10048 69176
rect 10100 69164 10106 69216
rect 1104 69114 10856 69136
rect 1104 69062 2582 69114
rect 2634 69062 2646 69114
rect 2698 69062 2710 69114
rect 2762 69062 2774 69114
rect 2826 69062 2838 69114
rect 2890 69062 5845 69114
rect 5897 69062 5909 69114
rect 5961 69062 5973 69114
rect 6025 69062 6037 69114
rect 6089 69062 6101 69114
rect 6153 69062 9109 69114
rect 9161 69062 9173 69114
rect 9225 69062 9237 69114
rect 9289 69062 9301 69114
rect 9353 69062 9365 69114
rect 9417 69062 10856 69114
rect 1104 69040 10856 69062
rect 3326 68960 3332 69012
rect 3384 69000 3390 69012
rect 6178 69000 6184 69012
rect 3384 68972 6184 69000
rect 3384 68960 3390 68972
rect 6178 68960 6184 68972
rect 6236 68960 6242 69012
rect 1394 68796 1400 68808
rect 1355 68768 1400 68796
rect 1394 68756 1400 68768
rect 1452 68756 1458 68808
rect 1486 68620 1492 68672
rect 1544 68660 1550 68672
rect 1581 68663 1639 68669
rect 1581 68660 1593 68663
rect 1544 68632 1593 68660
rect 1544 68620 1550 68632
rect 1581 68629 1593 68632
rect 1627 68629 1639 68663
rect 1581 68623 1639 68629
rect 1104 68570 10856 68592
rect 1104 68518 4213 68570
rect 4265 68518 4277 68570
rect 4329 68518 4341 68570
rect 4393 68518 4405 68570
rect 4457 68518 4469 68570
rect 4521 68518 7477 68570
rect 7529 68518 7541 68570
rect 7593 68518 7605 68570
rect 7657 68518 7669 68570
rect 7721 68518 7733 68570
rect 7785 68518 10856 68570
rect 1104 68496 10856 68518
rect 1394 68320 1400 68332
rect 1355 68292 1400 68320
rect 1394 68280 1400 68292
rect 1452 68280 1458 68332
rect 9858 68320 9864 68332
rect 9819 68292 9864 68320
rect 9858 68280 9864 68292
rect 9916 68280 9922 68332
rect 10042 68184 10048 68196
rect 10003 68156 10048 68184
rect 10042 68144 10048 68156
rect 10100 68144 10106 68196
rect 1581 68119 1639 68125
rect 1581 68085 1593 68119
rect 1627 68116 1639 68119
rect 1854 68116 1860 68128
rect 1627 68088 1860 68116
rect 1627 68085 1639 68088
rect 1581 68079 1639 68085
rect 1854 68076 1860 68088
rect 1912 68076 1918 68128
rect 1104 68026 10856 68048
rect 1104 67974 2582 68026
rect 2634 67974 2646 68026
rect 2698 67974 2710 68026
rect 2762 67974 2774 68026
rect 2826 67974 2838 68026
rect 2890 67974 5845 68026
rect 5897 67974 5909 68026
rect 5961 67974 5973 68026
rect 6025 67974 6037 68026
rect 6089 67974 6101 68026
rect 6153 67974 9109 68026
rect 9161 67974 9173 68026
rect 9225 67974 9237 68026
rect 9289 67974 9301 68026
rect 9353 67974 9365 68026
rect 9417 67974 10856 68026
rect 1104 67952 10856 67974
rect 1581 67915 1639 67921
rect 1581 67881 1593 67915
rect 1627 67912 1639 67915
rect 2130 67912 2136 67924
rect 1627 67884 2136 67912
rect 1627 67881 1639 67884
rect 1581 67875 1639 67881
rect 2130 67872 2136 67884
rect 2188 67872 2194 67924
rect 1946 67804 1952 67856
rect 2004 67844 2010 67856
rect 2041 67847 2099 67853
rect 2041 67844 2053 67847
rect 2004 67816 2053 67844
rect 2004 67804 2010 67816
rect 2041 67813 2053 67816
rect 2087 67813 2099 67847
rect 2041 67807 2099 67813
rect 1394 67708 1400 67720
rect 1355 67680 1400 67708
rect 1394 67668 1400 67680
rect 1452 67668 1458 67720
rect 2222 67708 2228 67720
rect 2183 67680 2228 67708
rect 2222 67668 2228 67680
rect 2280 67668 2286 67720
rect 9766 67668 9772 67720
rect 9824 67708 9830 67720
rect 9861 67711 9919 67717
rect 9861 67708 9873 67711
rect 9824 67680 9873 67708
rect 9824 67668 9830 67680
rect 9861 67677 9873 67680
rect 9907 67677 9919 67711
rect 9861 67671 9919 67677
rect 10042 67572 10048 67584
rect 10003 67544 10048 67572
rect 10042 67532 10048 67544
rect 10100 67532 10106 67584
rect 1104 67482 10856 67504
rect 1104 67430 4213 67482
rect 4265 67430 4277 67482
rect 4329 67430 4341 67482
rect 4393 67430 4405 67482
rect 4457 67430 4469 67482
rect 4521 67430 7477 67482
rect 7529 67430 7541 67482
rect 7593 67430 7605 67482
rect 7657 67430 7669 67482
rect 7721 67430 7733 67482
rect 7785 67430 10856 67482
rect 1104 67408 10856 67430
rect 1210 67192 1216 67244
rect 1268 67232 1274 67244
rect 1397 67235 1455 67241
rect 1397 67232 1409 67235
rect 1268 67204 1409 67232
rect 1268 67192 1274 67204
rect 1397 67201 1409 67204
rect 1443 67201 1455 67235
rect 2222 67232 2228 67244
rect 2183 67204 2228 67232
rect 1397 67195 1455 67201
rect 2222 67192 2228 67204
rect 2280 67192 2286 67244
rect 9582 67192 9588 67244
rect 9640 67232 9646 67244
rect 9861 67235 9919 67241
rect 9861 67232 9873 67235
rect 9640 67204 9873 67232
rect 9640 67192 9646 67204
rect 9861 67201 9873 67204
rect 9907 67201 9919 67235
rect 9861 67195 9919 67201
rect 2314 67124 2320 67176
rect 2372 67164 2378 67176
rect 3050 67164 3056 67176
rect 2372 67136 3056 67164
rect 2372 67124 2378 67136
rect 3050 67124 3056 67136
rect 3108 67124 3114 67176
rect 1578 67028 1584 67040
rect 1539 67000 1584 67028
rect 1578 66988 1584 67000
rect 1636 66988 1642 67040
rect 2041 67031 2099 67037
rect 2041 66997 2053 67031
rect 2087 67028 2099 67031
rect 2314 67028 2320 67040
rect 2087 67000 2320 67028
rect 2087 66997 2099 67000
rect 2041 66991 2099 66997
rect 2314 66988 2320 67000
rect 2372 66988 2378 67040
rect 3510 66988 3516 67040
rect 3568 67028 3574 67040
rect 4062 67028 4068 67040
rect 3568 67000 4068 67028
rect 3568 66988 3574 67000
rect 4062 66988 4068 67000
rect 4120 66988 4126 67040
rect 10042 67028 10048 67040
rect 10003 67000 10048 67028
rect 10042 66988 10048 67000
rect 10100 66988 10106 67040
rect 1104 66938 10856 66960
rect 1104 66886 2582 66938
rect 2634 66886 2646 66938
rect 2698 66886 2710 66938
rect 2762 66886 2774 66938
rect 2826 66886 2838 66938
rect 2890 66886 5845 66938
rect 5897 66886 5909 66938
rect 5961 66886 5973 66938
rect 6025 66886 6037 66938
rect 6089 66886 6101 66938
rect 6153 66886 9109 66938
rect 9161 66886 9173 66938
rect 9225 66886 9237 66938
rect 9289 66886 9301 66938
rect 9353 66886 9365 66938
rect 9417 66886 10856 66938
rect 1104 66864 10856 66886
rect 2961 66827 3019 66833
rect 2961 66793 2973 66827
rect 3007 66824 3019 66827
rect 9858 66824 9864 66836
rect 3007 66796 9864 66824
rect 3007 66793 3019 66796
rect 2961 66787 3019 66793
rect 9858 66784 9864 66796
rect 9916 66784 9922 66836
rect 2406 66716 2412 66768
rect 2464 66756 2470 66768
rect 2682 66756 2688 66768
rect 2464 66728 2688 66756
rect 2464 66716 2470 66728
rect 2682 66716 2688 66728
rect 2740 66716 2746 66768
rect 1302 66580 1308 66632
rect 1360 66620 1366 66632
rect 1397 66623 1455 66629
rect 1397 66620 1409 66623
rect 1360 66592 1409 66620
rect 1360 66580 1366 66592
rect 1397 66589 1409 66592
rect 1443 66589 1455 66623
rect 1397 66583 1455 66589
rect 2222 66580 2228 66632
rect 2280 66620 2286 66632
rect 2409 66623 2467 66629
rect 2409 66620 2421 66623
rect 2280 66592 2421 66620
rect 2280 66580 2286 66592
rect 2409 66589 2421 66592
rect 2455 66589 2467 66623
rect 2409 66583 2467 66589
rect 2498 66580 2504 66632
rect 2556 66620 2562 66632
rect 2685 66623 2743 66629
rect 2685 66620 2697 66623
rect 2556 66592 2697 66620
rect 2556 66580 2562 66592
rect 2685 66589 2697 66592
rect 2731 66589 2743 66623
rect 2685 66583 2743 66589
rect 2777 66623 2835 66629
rect 2777 66589 2789 66623
rect 2823 66620 2835 66623
rect 2866 66620 2872 66632
rect 2823 66592 2872 66620
rect 2823 66589 2835 66592
rect 2777 66583 2835 66589
rect 2866 66580 2872 66592
rect 2924 66580 2930 66632
rect 3510 66580 3516 66632
rect 3568 66620 3574 66632
rect 3786 66620 3792 66632
rect 3568 66592 3792 66620
rect 3568 66580 3574 66592
rect 3786 66580 3792 66592
rect 3844 66580 3850 66632
rect 2593 66555 2651 66561
rect 2593 66521 2605 66555
rect 2639 66521 2651 66555
rect 2593 66515 2651 66521
rect 1581 66487 1639 66493
rect 1581 66453 1593 66487
rect 1627 66484 1639 66487
rect 2406 66484 2412 66496
rect 1627 66456 2412 66484
rect 1627 66453 1639 66456
rect 1581 66447 1639 66453
rect 2406 66444 2412 66456
rect 2464 66444 2470 66496
rect 2608 66484 2636 66515
rect 2608 66456 10916 66484
rect 1104 66394 10856 66416
rect 1104 66342 4213 66394
rect 4265 66342 4277 66394
rect 4329 66342 4341 66394
rect 4393 66342 4405 66394
rect 4457 66342 4469 66394
rect 4521 66342 7477 66394
rect 7529 66342 7541 66394
rect 7593 66342 7605 66394
rect 7657 66342 7669 66394
rect 7721 66342 7733 66394
rect 7785 66342 10856 66394
rect 1104 66320 10856 66342
rect 2222 66280 2228 66292
rect 1412 66252 2228 66280
rect 1412 66153 1440 66252
rect 2222 66240 2228 66252
rect 2280 66280 2286 66292
rect 2280 66252 2820 66280
rect 2280 66240 2286 66252
rect 1670 66212 1676 66224
rect 1631 66184 1676 66212
rect 1670 66172 1676 66184
rect 1728 66172 1734 66224
rect 1397 66147 1455 66153
rect 1397 66113 1409 66147
rect 1443 66113 1455 66147
rect 1397 66107 1455 66113
rect 1581 66147 1639 66153
rect 1581 66113 1593 66147
rect 1627 66113 1639 66147
rect 1581 66107 1639 66113
rect 1765 66147 1823 66153
rect 1765 66113 1777 66147
rect 1811 66113 1823 66147
rect 2332 66144 2360 66252
rect 2792 66212 2820 66252
rect 2866 66240 2872 66292
rect 2924 66280 2930 66292
rect 10888 66289 10916 66456
rect 10873 66283 10931 66289
rect 2924 66252 3832 66280
rect 2924 66240 2930 66252
rect 3694 66212 3700 66224
rect 2792 66184 3464 66212
rect 3655 66184 3700 66212
rect 2409 66147 2467 66153
rect 2409 66144 2421 66147
rect 2332 66116 2421 66144
rect 1765 66107 1823 66113
rect 2409 66113 2421 66116
rect 2455 66113 2467 66147
rect 2409 66107 2467 66113
rect 750 66036 756 66088
rect 808 66076 814 66088
rect 1596 66076 1624 66107
rect 808 66048 1624 66076
rect 1780 66076 1808 66107
rect 2498 66104 2504 66156
rect 2556 66153 2562 66156
rect 2556 66147 2605 66153
rect 2556 66113 2559 66147
rect 2593 66113 2605 66147
rect 2682 66144 2688 66156
rect 2643 66116 2688 66144
rect 2556 66107 2605 66113
rect 2556 66104 2562 66107
rect 2682 66104 2688 66116
rect 2740 66104 2746 66156
rect 2777 66147 2835 66153
rect 2777 66113 2789 66147
rect 2823 66144 2835 66147
rect 2866 66144 2872 66156
rect 2823 66116 2872 66144
rect 2823 66113 2835 66116
rect 2777 66107 2835 66113
rect 2792 66076 2820 66107
rect 2866 66104 2872 66116
rect 2924 66104 2930 66156
rect 3436 66153 3464 66184
rect 3694 66172 3700 66184
rect 3752 66172 3758 66224
rect 3421 66147 3479 66153
rect 3421 66113 3433 66147
rect 3467 66113 3479 66147
rect 3602 66144 3608 66156
rect 3563 66116 3608 66144
rect 3421 66107 3479 66113
rect 3602 66104 3608 66116
rect 3660 66104 3666 66156
rect 3804 66153 3832 66252
rect 10873 66249 10885 66283
rect 10919 66249 10931 66283
rect 10873 66243 10931 66249
rect 9769 66215 9827 66221
rect 9769 66181 9781 66215
rect 9815 66212 9827 66215
rect 11057 66215 11115 66221
rect 11057 66212 11069 66215
rect 9815 66184 11069 66212
rect 9815 66181 9827 66184
rect 9769 66175 9827 66181
rect 11057 66181 11069 66184
rect 11103 66181 11115 66215
rect 11057 66175 11115 66181
rect 3789 66147 3847 66153
rect 3789 66113 3801 66147
rect 3835 66144 3847 66147
rect 3970 66144 3976 66156
rect 3835 66116 3976 66144
rect 3835 66113 3847 66116
rect 3789 66107 3847 66113
rect 3970 66104 3976 66116
rect 4028 66104 4034 66156
rect 9674 66104 9680 66156
rect 9732 66144 9738 66156
rect 9861 66147 9919 66153
rect 9861 66144 9873 66147
rect 9732 66116 9873 66144
rect 9732 66104 9738 66116
rect 9861 66113 9873 66116
rect 9907 66113 9919 66147
rect 9861 66107 9919 66113
rect 9766 66076 9772 66088
rect 1780 66048 2820 66076
rect 2976 66048 9772 66076
rect 808 66036 814 66048
rect 2976 66017 3004 66048
rect 9766 66036 9772 66048
rect 9824 66036 9830 66088
rect 2961 66011 3019 66017
rect 2961 65977 2973 66011
rect 3007 65977 3019 66011
rect 2961 65971 3019 65977
rect 3973 66011 4031 66017
rect 3973 65977 3985 66011
rect 4019 66008 4031 66011
rect 10965 66011 11023 66017
rect 10965 66008 10977 66011
rect 4019 65980 10977 66008
rect 4019 65977 4031 65980
rect 3973 65971 4031 65977
rect 10965 65977 10977 65980
rect 11011 65977 11023 66011
rect 10965 65971 11023 65977
rect 1949 65943 2007 65949
rect 1949 65909 1961 65943
rect 1995 65940 2007 65943
rect 9769 65943 9827 65949
rect 9769 65940 9781 65943
rect 1995 65912 9781 65940
rect 1995 65909 2007 65912
rect 1949 65903 2007 65909
rect 9769 65909 9781 65912
rect 9815 65909 9827 65943
rect 10042 65940 10048 65952
rect 10003 65912 10048 65940
rect 9769 65903 9827 65909
rect 10042 65900 10048 65912
rect 10100 65900 10106 65952
rect 1104 65850 10856 65872
rect 1104 65798 2582 65850
rect 2634 65798 2646 65850
rect 2698 65798 2710 65850
rect 2762 65798 2774 65850
rect 2826 65798 2838 65850
rect 2890 65798 5845 65850
rect 5897 65798 5909 65850
rect 5961 65798 5973 65850
rect 6025 65798 6037 65850
rect 6089 65798 6101 65850
rect 6153 65798 9109 65850
rect 9161 65798 9173 65850
rect 9225 65798 9237 65850
rect 9289 65798 9301 65850
rect 9353 65798 9365 65850
rect 9417 65798 10856 65850
rect 1104 65776 10856 65798
rect 3602 65736 3608 65748
rect 1136 65708 3608 65736
rect 1026 65356 1032 65408
rect 1084 65396 1090 65408
rect 1136 65396 1164 65708
rect 3602 65696 3608 65708
rect 3660 65696 3666 65748
rect 3786 65668 3792 65680
rect 3252 65640 3792 65668
rect 3252 65612 3280 65640
rect 3786 65628 3792 65640
rect 3844 65628 3850 65680
rect 2222 65560 2228 65612
rect 2280 65600 2286 65612
rect 2961 65603 3019 65609
rect 2961 65600 2973 65603
rect 2280 65572 2973 65600
rect 2280 65560 2286 65572
rect 2961 65569 2973 65572
rect 3007 65569 3019 65603
rect 2961 65563 3019 65569
rect 3234 65560 3240 65612
rect 3292 65600 3298 65612
rect 3292 65572 3385 65600
rect 3292 65560 3298 65572
rect 3970 65560 3976 65612
rect 4028 65600 4034 65612
rect 4065 65603 4123 65609
rect 4065 65600 4077 65603
rect 4028 65572 4077 65600
rect 4028 65560 4034 65572
rect 4065 65569 4077 65572
rect 4111 65569 4123 65603
rect 4065 65563 4123 65569
rect 1394 65532 1400 65544
rect 1355 65504 1400 65532
rect 1394 65492 1400 65504
rect 1452 65492 1458 65544
rect 3510 65492 3516 65544
rect 3568 65532 3574 65544
rect 3789 65535 3847 65541
rect 3789 65532 3801 65535
rect 3568 65504 3801 65532
rect 3568 65492 3574 65504
rect 3789 65501 3801 65504
rect 3835 65501 3847 65535
rect 9858 65532 9864 65544
rect 9819 65504 9864 65532
rect 3789 65495 3847 65501
rect 9858 65492 9864 65504
rect 9916 65492 9922 65544
rect 1084 65368 1164 65396
rect 1581 65399 1639 65405
rect 1084 65356 1090 65368
rect 1581 65365 1593 65399
rect 1627 65396 1639 65399
rect 1670 65396 1676 65408
rect 1627 65368 1676 65396
rect 1627 65365 1639 65368
rect 1581 65359 1639 65365
rect 1670 65356 1676 65368
rect 1728 65356 1734 65408
rect 10042 65396 10048 65408
rect 10003 65368 10048 65396
rect 10042 65356 10048 65368
rect 10100 65356 10106 65408
rect 1104 65306 10856 65328
rect 1104 65254 4213 65306
rect 4265 65254 4277 65306
rect 4329 65254 4341 65306
rect 4393 65254 4405 65306
rect 4457 65254 4469 65306
rect 4521 65254 7477 65306
rect 7529 65254 7541 65306
rect 7593 65254 7605 65306
rect 7657 65254 7669 65306
rect 7721 65254 7733 65306
rect 7785 65254 10856 65306
rect 1104 65232 10856 65254
rect 842 65152 848 65204
rect 900 65192 906 65204
rect 1210 65192 1216 65204
rect 900 65164 1216 65192
rect 900 65152 906 65164
rect 1210 65152 1216 65164
rect 1268 65152 1274 65204
rect 2961 65195 3019 65201
rect 2961 65161 2973 65195
rect 3007 65192 3019 65195
rect 9582 65192 9588 65204
rect 3007 65164 9588 65192
rect 3007 65161 3019 65164
rect 2961 65155 3019 65161
rect 9582 65152 9588 65164
rect 9640 65152 9646 65204
rect 2038 65084 2044 65136
rect 2096 65124 2102 65136
rect 2593 65127 2651 65133
rect 2096 65096 2544 65124
rect 2096 65084 2102 65096
rect 1302 65016 1308 65068
rect 1360 65056 1366 65068
rect 1397 65059 1455 65065
rect 1397 65056 1409 65059
rect 1360 65028 1409 65056
rect 1360 65016 1366 65028
rect 1397 65025 1409 65028
rect 1443 65025 1455 65059
rect 1397 65019 1455 65025
rect 2222 65016 2228 65068
rect 2280 65056 2286 65068
rect 2409 65059 2467 65065
rect 2409 65056 2421 65059
rect 2280 65028 2421 65056
rect 2280 65016 2286 65028
rect 2409 65025 2421 65028
rect 2455 65025 2467 65059
rect 2516 65056 2544 65096
rect 2593 65093 2605 65127
rect 2639 65124 2651 65127
rect 5350 65124 5356 65136
rect 2639 65096 5356 65124
rect 2639 65093 2651 65096
rect 2593 65087 2651 65093
rect 5350 65084 5356 65096
rect 5408 65084 5414 65136
rect 2685 65059 2743 65065
rect 2685 65056 2697 65059
rect 2516 65028 2697 65056
rect 2409 65019 2467 65025
rect 2685 65025 2697 65028
rect 2731 65025 2743 65059
rect 2685 65019 2743 65025
rect 2777 65059 2835 65065
rect 2777 65025 2789 65059
rect 2823 65056 2835 65059
rect 2958 65056 2964 65068
rect 2823 65028 2964 65056
rect 2823 65025 2835 65028
rect 2777 65019 2835 65025
rect 2958 65016 2964 65028
rect 3016 65016 3022 65068
rect 2498 64948 2504 65000
rect 2556 64988 2562 65000
rect 6638 64988 6644 65000
rect 2556 64960 6644 64988
rect 2556 64948 2562 64960
rect 6638 64948 6644 64960
rect 6696 64948 6702 65000
rect 1581 64923 1639 64929
rect 1581 64889 1593 64923
rect 1627 64920 1639 64923
rect 2222 64920 2228 64932
rect 1627 64892 2228 64920
rect 1627 64889 1639 64892
rect 1581 64883 1639 64889
rect 2222 64880 2228 64892
rect 2280 64880 2286 64932
rect 1104 64762 10856 64784
rect 1104 64710 2582 64762
rect 2634 64710 2646 64762
rect 2698 64710 2710 64762
rect 2762 64710 2774 64762
rect 2826 64710 2838 64762
rect 2890 64710 5845 64762
rect 5897 64710 5909 64762
rect 5961 64710 5973 64762
rect 6025 64710 6037 64762
rect 6089 64710 6101 64762
rect 6153 64710 9109 64762
rect 9161 64710 9173 64762
rect 9225 64710 9237 64762
rect 9289 64710 9301 64762
rect 9353 64710 9365 64762
rect 9417 64710 10856 64762
rect 1104 64688 10856 64710
rect 937 64651 995 64657
rect 937 64617 949 64651
rect 983 64648 995 64651
rect 2501 64651 2559 64657
rect 2501 64648 2513 64651
rect 983 64620 2513 64648
rect 983 64617 995 64620
rect 937 64611 995 64617
rect 2501 64617 2513 64620
rect 2547 64617 2559 64651
rect 2501 64611 2559 64617
rect 2041 64583 2099 64589
rect 2041 64549 2053 64583
rect 2087 64580 2099 64583
rect 9858 64580 9864 64592
rect 2087 64552 9864 64580
rect 2087 64549 2099 64552
rect 2041 64543 2099 64549
rect 9858 64540 9864 64552
rect 9916 64540 9922 64592
rect 2958 64512 2964 64524
rect 1872 64484 2964 64512
rect 1394 64404 1400 64456
rect 1452 64444 1458 64456
rect 1489 64447 1547 64453
rect 1489 64444 1501 64447
rect 1452 64416 1501 64444
rect 1452 64404 1458 64416
rect 1489 64413 1501 64416
rect 1535 64413 1547 64447
rect 1762 64444 1768 64456
rect 1723 64416 1768 64444
rect 1489 64407 1547 64413
rect 1762 64404 1768 64416
rect 1820 64404 1826 64456
rect 1872 64453 1900 64484
rect 2958 64472 2964 64484
rect 3016 64472 3022 64524
rect 1857 64447 1915 64453
rect 1857 64413 1869 64447
rect 1903 64413 1915 64447
rect 1857 64407 1915 64413
rect 2685 64447 2743 64453
rect 2685 64413 2697 64447
rect 2731 64444 2743 64447
rect 2774 64444 2780 64456
rect 2731 64416 2780 64444
rect 2731 64413 2743 64416
rect 2685 64407 2743 64413
rect 2774 64404 2780 64416
rect 2832 64404 2838 64456
rect 2866 64404 2872 64456
rect 2924 64444 2930 64456
rect 3050 64444 3056 64456
rect 2924 64416 3056 64444
rect 2924 64404 2930 64416
rect 3050 64404 3056 64416
rect 3108 64404 3114 64456
rect 9766 64404 9772 64456
rect 9824 64444 9830 64456
rect 9861 64447 9919 64453
rect 9861 64444 9873 64447
rect 9824 64416 9873 64444
rect 9824 64404 9830 64416
rect 9861 64413 9873 64416
rect 9907 64413 9919 64447
rect 9861 64407 9919 64413
rect 1673 64379 1731 64385
rect 1673 64345 1685 64379
rect 1719 64345 1731 64379
rect 7190 64376 7196 64388
rect 1673 64339 1731 64345
rect 1964 64348 7196 64376
rect 1688 64308 1716 64339
rect 1964 64308 1992 64348
rect 7190 64336 7196 64348
rect 7248 64336 7254 64388
rect 10042 64308 10048 64320
rect 1688 64280 1992 64308
rect 10003 64280 10048 64308
rect 10042 64268 10048 64280
rect 10100 64268 10106 64320
rect 1104 64218 10856 64240
rect 1104 64166 4213 64218
rect 4265 64166 4277 64218
rect 4329 64166 4341 64218
rect 4393 64166 4405 64218
rect 4457 64166 4469 64218
rect 4521 64166 7477 64218
rect 7529 64166 7541 64218
rect 7593 64166 7605 64218
rect 7657 64166 7669 64218
rect 7721 64166 7733 64218
rect 7785 64166 10856 64218
rect 1104 64144 10856 64166
rect 1486 64064 1492 64116
rect 1544 64104 1550 64116
rect 3053 64107 3111 64113
rect 1544 64076 1716 64104
rect 1544 64064 1550 64076
rect 1688 64036 1716 64076
rect 3053 64073 3065 64107
rect 3099 64104 3111 64107
rect 9674 64104 9680 64116
rect 3099 64076 9680 64104
rect 3099 64073 3111 64076
rect 3053 64067 3111 64073
rect 9674 64064 9680 64076
rect 9732 64064 9738 64116
rect 1765 64039 1823 64045
rect 1765 64036 1777 64039
rect 1688 64008 1777 64036
rect 1765 64005 1777 64008
rect 1811 64005 1823 64039
rect 1765 63999 1823 64005
rect 2685 64039 2743 64045
rect 2685 64005 2697 64039
rect 2731 64036 2743 64039
rect 8386 64036 8392 64048
rect 2731 64008 8392 64036
rect 2731 64005 2743 64008
rect 2685 63999 2743 64005
rect 8386 63996 8392 64008
rect 8444 63996 8450 64048
rect 1486 63968 1492 63980
rect 1447 63940 1492 63968
rect 1486 63928 1492 63940
rect 1544 63928 1550 63980
rect 1673 63971 1731 63977
rect 1673 63937 1685 63971
rect 1719 63937 1731 63971
rect 1673 63931 1731 63937
rect 1903 63971 1961 63977
rect 1903 63937 1915 63971
rect 1949 63968 1961 63971
rect 2498 63968 2504 63980
rect 1949 63940 2084 63968
rect 2459 63940 2504 63968
rect 1949 63937 1961 63940
rect 1903 63931 1961 63937
rect 1688 63764 1716 63931
rect 2056 63900 2084 63940
rect 2498 63928 2504 63940
rect 2556 63928 2562 63980
rect 2774 63968 2780 63980
rect 2735 63940 2780 63968
rect 2774 63928 2780 63940
rect 2832 63928 2838 63980
rect 2869 63971 2927 63977
rect 2869 63937 2881 63971
rect 2915 63968 2927 63971
rect 2958 63968 2964 63980
rect 2915 63940 2964 63968
rect 2915 63937 2927 63940
rect 2869 63931 2927 63937
rect 2884 63900 2912 63931
rect 2958 63928 2964 63940
rect 3016 63928 3022 63980
rect 9858 63968 9864 63980
rect 9819 63940 9864 63968
rect 9858 63928 9864 63940
rect 9916 63928 9922 63980
rect 2056 63872 2912 63900
rect 2041 63835 2099 63841
rect 2041 63801 2053 63835
rect 2087 63832 2099 63835
rect 9766 63832 9772 63844
rect 2087 63804 9772 63832
rect 2087 63801 2099 63804
rect 2041 63795 2099 63801
rect 9766 63792 9772 63804
rect 9824 63792 9830 63844
rect 8294 63764 8300 63776
rect 1688 63736 8300 63764
rect 8294 63724 8300 63736
rect 8352 63724 8358 63776
rect 10042 63764 10048 63776
rect 10003 63736 10048 63764
rect 10042 63724 10048 63736
rect 10100 63724 10106 63776
rect 1104 63674 10856 63696
rect 1104 63622 2582 63674
rect 2634 63622 2646 63674
rect 2698 63622 2710 63674
rect 2762 63622 2774 63674
rect 2826 63622 2838 63674
rect 2890 63622 5845 63674
rect 5897 63622 5909 63674
rect 5961 63622 5973 63674
rect 6025 63622 6037 63674
rect 6089 63622 6101 63674
rect 6153 63622 9109 63674
rect 9161 63622 9173 63674
rect 9225 63622 9237 63674
rect 9289 63622 9301 63674
rect 9353 63622 9365 63674
rect 9417 63622 10856 63674
rect 1104 63600 10856 63622
rect 1762 63520 1768 63572
rect 1820 63560 1826 63572
rect 2038 63560 2044 63572
rect 1820 63532 2044 63560
rect 1820 63520 1826 63532
rect 2038 63520 2044 63532
rect 2096 63520 2102 63572
rect 2314 63520 2320 63572
rect 2372 63560 2378 63572
rect 2498 63560 2504 63572
rect 2372 63532 2504 63560
rect 2372 63520 2378 63532
rect 2498 63520 2504 63532
rect 2556 63520 2562 63572
rect 2133 63495 2191 63501
rect 2133 63461 2145 63495
rect 2179 63492 2191 63495
rect 9858 63492 9864 63504
rect 2179 63464 9864 63492
rect 2179 63461 2191 63464
rect 2133 63455 2191 63461
rect 9858 63452 9864 63464
rect 9916 63452 9922 63504
rect 2866 63384 2872 63436
rect 2924 63424 2930 63436
rect 3326 63424 3332 63436
rect 2924 63396 3332 63424
rect 2924 63384 2930 63396
rect 3326 63384 3332 63396
rect 3384 63424 3390 63436
rect 3510 63424 3516 63436
rect 3384 63396 3516 63424
rect 3384 63384 3390 63396
rect 3510 63384 3516 63396
rect 3568 63384 3574 63436
rect 1486 63316 1492 63368
rect 1544 63356 1550 63368
rect 1581 63359 1639 63365
rect 1581 63356 1593 63359
rect 1544 63328 1593 63356
rect 1544 63316 1550 63328
rect 1581 63325 1593 63328
rect 1627 63325 1639 63359
rect 1854 63356 1860 63368
rect 1815 63328 1860 63356
rect 1581 63319 1639 63325
rect 1854 63316 1860 63328
rect 1912 63316 1918 63368
rect 1949 63359 2007 63365
rect 1949 63325 1961 63359
rect 1995 63356 2007 63359
rect 2038 63356 2044 63368
rect 1995 63328 2044 63356
rect 1995 63325 2007 63328
rect 1949 63319 2007 63325
rect 2038 63316 2044 63328
rect 2096 63316 2102 63368
rect 2774 63316 2780 63368
rect 2832 63356 2838 63368
rect 3970 63356 3976 63368
rect 2832 63328 2877 63356
rect 3931 63328 3976 63356
rect 2832 63316 2838 63328
rect 3970 63316 3976 63328
rect 4028 63316 4034 63368
rect 9858 63356 9864 63368
rect 9819 63328 9864 63356
rect 9858 63316 9864 63328
rect 9916 63316 9922 63368
rect 1765 63291 1823 63297
rect 1765 63257 1777 63291
rect 1811 63257 1823 63291
rect 6914 63288 6920 63300
rect 1765 63251 1823 63257
rect 2056 63260 6920 63288
rect 1780 63220 1808 63251
rect 2056 63220 2084 63260
rect 6914 63248 6920 63260
rect 6972 63248 6978 63300
rect 2590 63220 2596 63232
rect 1780 63192 2084 63220
rect 2551 63192 2596 63220
rect 2590 63180 2596 63192
rect 2648 63180 2654 63232
rect 2682 63180 2688 63232
rect 2740 63220 2746 63232
rect 3789 63223 3847 63229
rect 3789 63220 3801 63223
rect 2740 63192 3801 63220
rect 2740 63180 2746 63192
rect 3789 63189 3801 63192
rect 3835 63189 3847 63223
rect 10042 63220 10048 63232
rect 10003 63192 10048 63220
rect 3789 63183 3847 63189
rect 10042 63180 10048 63192
rect 10100 63180 10106 63232
rect 1104 63130 10856 63152
rect 1104 63078 4213 63130
rect 4265 63078 4277 63130
rect 4329 63078 4341 63130
rect 4393 63078 4405 63130
rect 4457 63078 4469 63130
rect 4521 63078 7477 63130
rect 7529 63078 7541 63130
rect 7593 63078 7605 63130
rect 7657 63078 7669 63130
rect 7721 63078 7733 63130
rect 7785 63078 10856 63130
rect 1104 63056 10856 63078
rect 2685 63019 2743 63025
rect 2685 62985 2697 63019
rect 2731 63016 2743 63019
rect 2958 63016 2964 63028
rect 2731 62988 2964 63016
rect 2731 62985 2743 62988
rect 2685 62979 2743 62985
rect 2958 62976 2964 62988
rect 3016 63016 3022 63028
rect 3016 62988 3096 63016
rect 3016 62976 3022 62988
rect 1857 62951 1915 62957
rect 1857 62917 1869 62951
rect 1903 62948 1915 62951
rect 1903 62920 3004 62948
rect 1903 62917 1915 62920
rect 1857 62911 1915 62917
rect 1486 62840 1492 62892
rect 1544 62880 1550 62892
rect 1673 62883 1731 62889
rect 1673 62880 1685 62883
rect 1544 62852 1685 62880
rect 1544 62840 1550 62852
rect 1673 62849 1685 62852
rect 1719 62880 1731 62883
rect 1762 62880 1768 62892
rect 1719 62852 1768 62880
rect 1719 62849 1731 62852
rect 1673 62843 1731 62849
rect 1762 62840 1768 62852
rect 1820 62840 1826 62892
rect 1946 62880 1952 62892
rect 1907 62852 1952 62880
rect 1946 62840 1952 62852
rect 2004 62840 2010 62892
rect 2038 62840 2044 62892
rect 2096 62880 2102 62892
rect 2685 62883 2743 62889
rect 2685 62880 2697 62883
rect 2096 62852 2697 62880
rect 2096 62840 2102 62852
rect 2685 62849 2697 62852
rect 2731 62849 2743 62883
rect 2685 62843 2743 62849
rect 2777 62883 2835 62889
rect 2777 62849 2789 62883
rect 2823 62880 2835 62883
rect 2866 62880 2872 62892
rect 2823 62852 2872 62880
rect 2823 62849 2835 62852
rect 2777 62843 2835 62849
rect 2866 62840 2872 62852
rect 2924 62840 2930 62892
rect 2590 62812 2596 62824
rect 1964 62784 2596 62812
rect 1964 62756 1992 62784
rect 2590 62772 2596 62784
rect 2648 62772 2654 62824
rect 1946 62704 1952 62756
rect 2004 62704 2010 62756
rect 2038 62704 2044 62756
rect 2096 62744 2102 62756
rect 2682 62744 2688 62756
rect 2096 62716 2688 62744
rect 2096 62704 2102 62716
rect 2682 62704 2688 62716
rect 2740 62704 2746 62756
rect 2976 62744 3004 62920
rect 3068 62889 3096 62988
rect 3053 62883 3111 62889
rect 3053 62849 3065 62883
rect 3099 62849 3111 62883
rect 3053 62843 3111 62849
rect 8478 62744 8484 62756
rect 2976 62716 8484 62744
rect 8478 62704 8484 62716
rect 8536 62704 8542 62756
rect 2225 62679 2283 62685
rect 2225 62645 2237 62679
rect 2271 62676 2283 62679
rect 9858 62676 9864 62688
rect 2271 62648 9864 62676
rect 2271 62645 2283 62648
rect 2225 62639 2283 62645
rect 9858 62636 9864 62648
rect 9916 62636 9922 62688
rect 1104 62586 10856 62608
rect 1104 62534 2582 62586
rect 2634 62534 2646 62586
rect 2698 62534 2710 62586
rect 2762 62534 2774 62586
rect 2826 62534 2838 62586
rect 2890 62534 5845 62586
rect 5897 62534 5909 62586
rect 5961 62534 5973 62586
rect 6025 62534 6037 62586
rect 6089 62534 6101 62586
rect 6153 62534 9109 62586
rect 9161 62534 9173 62586
rect 9225 62534 9237 62586
rect 9289 62534 9301 62586
rect 9353 62534 9365 62586
rect 9417 62534 10856 62586
rect 1104 62512 10856 62534
rect 2038 62432 2044 62484
rect 2096 62472 2102 62484
rect 2406 62472 2412 62484
rect 2096 62444 2412 62472
rect 2096 62432 2102 62444
rect 2406 62432 2412 62444
rect 2464 62432 2470 62484
rect 1762 62296 1768 62348
rect 1820 62336 1826 62348
rect 2961 62339 3019 62345
rect 2961 62336 2973 62339
rect 1820 62308 2973 62336
rect 1820 62296 1826 62308
rect 2961 62305 2973 62308
rect 3007 62305 3019 62339
rect 3234 62336 3240 62348
rect 3195 62308 3240 62336
rect 2961 62299 3019 62305
rect 3234 62296 3240 62308
rect 3292 62296 3298 62348
rect 1673 62271 1731 62277
rect 1673 62237 1685 62271
rect 1719 62268 1731 62271
rect 9861 62271 9919 62277
rect 1719 62240 2774 62268
rect 1719 62237 1731 62240
rect 1673 62231 1731 62237
rect 2746 62200 2774 62240
rect 9861 62237 9873 62271
rect 9907 62268 9919 62271
rect 11425 62271 11483 62277
rect 11425 62268 11437 62271
rect 9907 62240 11437 62268
rect 9907 62237 9919 62240
rect 9861 62231 9919 62237
rect 11425 62237 11437 62240
rect 11471 62237 11483 62271
rect 11425 62231 11483 62237
rect 3786 62200 3792 62212
rect 2746 62172 3792 62200
rect 3786 62160 3792 62172
rect 3844 62160 3850 62212
rect 1486 62132 1492 62144
rect 1447 62104 1492 62132
rect 1486 62092 1492 62104
rect 1544 62092 1550 62144
rect 1946 62092 1952 62144
rect 2004 62132 2010 62144
rect 2130 62132 2136 62144
rect 2004 62104 2136 62132
rect 2004 62092 2010 62104
rect 2130 62092 2136 62104
rect 2188 62092 2194 62144
rect 10042 62132 10048 62144
rect 10003 62104 10048 62132
rect 10042 62092 10048 62104
rect 10100 62092 10106 62144
rect 1104 62042 10856 62064
rect 1104 61990 4213 62042
rect 4265 61990 4277 62042
rect 4329 61990 4341 62042
rect 4393 61990 4405 62042
rect 4457 61990 4469 62042
rect 4521 61990 7477 62042
rect 7529 61990 7541 62042
rect 7593 61990 7605 62042
rect 7657 61990 7669 62042
rect 7721 61990 7733 62042
rect 7785 61990 10856 62042
rect 1104 61968 10856 61990
rect 1673 61795 1731 61801
rect 1673 61761 1685 61795
rect 1719 61761 1731 61795
rect 2314 61792 2320 61804
rect 2275 61764 2320 61792
rect 1673 61755 1731 61761
rect 1688 61724 1716 61755
rect 2314 61752 2320 61764
rect 2372 61752 2378 61804
rect 9861 61795 9919 61801
rect 9861 61761 9873 61795
rect 9907 61792 9919 61795
rect 11241 61795 11299 61801
rect 11241 61792 11253 61795
rect 9907 61764 11253 61792
rect 9907 61761 9919 61764
rect 9861 61755 9919 61761
rect 11241 61761 11253 61764
rect 11287 61761 11299 61795
rect 11241 61755 11299 61761
rect 3694 61724 3700 61736
rect 1688 61696 3700 61724
rect 3694 61684 3700 61696
rect 3752 61684 3758 61736
rect 1394 61548 1400 61600
rect 1452 61588 1458 61600
rect 1489 61591 1547 61597
rect 1489 61588 1501 61591
rect 1452 61560 1501 61588
rect 1452 61548 1458 61560
rect 1489 61557 1501 61560
rect 1535 61557 1547 61591
rect 1489 61551 1547 61557
rect 1762 61548 1768 61600
rect 1820 61588 1826 61600
rect 2133 61591 2191 61597
rect 2133 61588 2145 61591
rect 1820 61560 2145 61588
rect 1820 61548 1826 61560
rect 2133 61557 2145 61560
rect 2179 61557 2191 61591
rect 10042 61588 10048 61600
rect 10003 61560 10048 61588
rect 2133 61551 2191 61557
rect 10042 61548 10048 61560
rect 10100 61548 10106 61600
rect 1104 61498 10856 61520
rect 1104 61446 2582 61498
rect 2634 61446 2646 61498
rect 2698 61446 2710 61498
rect 2762 61446 2774 61498
rect 2826 61446 2838 61498
rect 2890 61446 5845 61498
rect 5897 61446 5909 61498
rect 5961 61446 5973 61498
rect 6025 61446 6037 61498
rect 6089 61446 6101 61498
rect 6153 61446 9109 61498
rect 9161 61446 9173 61498
rect 9225 61446 9237 61498
rect 9289 61446 9301 61498
rect 9353 61446 9365 61498
rect 9417 61446 10856 61498
rect 1104 61424 10856 61446
rect 1673 61183 1731 61189
rect 1673 61149 1685 61183
rect 1719 61180 1731 61183
rect 2314 61180 2320 61192
rect 1719 61152 2320 61180
rect 1719 61149 1731 61152
rect 1673 61143 1731 61149
rect 2314 61140 2320 61152
rect 2372 61140 2378 61192
rect 1486 61044 1492 61056
rect 1447 61016 1492 61044
rect 1486 61004 1492 61016
rect 1544 61004 1550 61056
rect 1104 60954 10856 60976
rect 1104 60902 4213 60954
rect 4265 60902 4277 60954
rect 4329 60902 4341 60954
rect 4393 60902 4405 60954
rect 4457 60902 4469 60954
rect 4521 60902 7477 60954
rect 7529 60902 7541 60954
rect 7593 60902 7605 60954
rect 7657 60902 7669 60954
rect 7721 60902 7733 60954
rect 7785 60902 10856 60954
rect 1104 60880 10856 60902
rect 1673 60707 1731 60713
rect 1673 60673 1685 60707
rect 1719 60704 1731 60707
rect 9861 60707 9919 60713
rect 1719 60676 2774 60704
rect 1719 60673 1731 60676
rect 1673 60667 1731 60673
rect 2746 60636 2774 60676
rect 9861 60673 9873 60707
rect 9907 60704 9919 60707
rect 11057 60707 11115 60713
rect 11057 60704 11069 60707
rect 9907 60676 11069 60704
rect 9907 60673 9919 60676
rect 9861 60667 9919 60673
rect 11057 60673 11069 60676
rect 11103 60673 11115 60707
rect 11057 60667 11115 60673
rect 3234 60636 3240 60648
rect 2746 60608 3240 60636
rect 3234 60596 3240 60608
rect 3292 60596 3298 60648
rect 10042 60568 10048 60580
rect 10003 60540 10048 60568
rect 10042 60528 10048 60540
rect 10100 60528 10106 60580
rect 1394 60460 1400 60512
rect 1452 60500 1458 60512
rect 1489 60503 1547 60509
rect 1489 60500 1501 60503
rect 1452 60472 1501 60500
rect 1452 60460 1458 60472
rect 1489 60469 1501 60472
rect 1535 60469 1547 60503
rect 1489 60463 1547 60469
rect 1104 60410 10856 60432
rect 1104 60358 2582 60410
rect 2634 60358 2646 60410
rect 2698 60358 2710 60410
rect 2762 60358 2774 60410
rect 2826 60358 2838 60410
rect 2890 60358 5845 60410
rect 5897 60358 5909 60410
rect 5961 60358 5973 60410
rect 6025 60358 6037 60410
rect 6089 60358 6101 60410
rect 6153 60358 9109 60410
rect 9161 60358 9173 60410
rect 9225 60358 9237 60410
rect 9289 60358 9301 60410
rect 9353 60358 9365 60410
rect 9417 60358 10856 60410
rect 1104 60336 10856 60358
rect 1673 60095 1731 60101
rect 1673 60061 1685 60095
rect 1719 60092 1731 60095
rect 3418 60092 3424 60104
rect 1719 60064 3424 60092
rect 1719 60061 1731 60064
rect 1673 60055 1731 60061
rect 3418 60052 3424 60064
rect 3476 60052 3482 60104
rect 9766 60052 9772 60104
rect 9824 60092 9830 60104
rect 9861 60095 9919 60101
rect 9861 60092 9873 60095
rect 9824 60064 9873 60092
rect 9824 60052 9830 60064
rect 9861 60061 9873 60064
rect 9907 60061 9919 60095
rect 9861 60055 9919 60061
rect 1486 59956 1492 59968
rect 1447 59928 1492 59956
rect 1486 59916 1492 59928
rect 1544 59916 1550 59968
rect 10042 59956 10048 59968
rect 10003 59928 10048 59956
rect 10042 59916 10048 59928
rect 10100 59916 10106 59968
rect 1104 59866 10856 59888
rect 1104 59814 4213 59866
rect 4265 59814 4277 59866
rect 4329 59814 4341 59866
rect 4393 59814 4405 59866
rect 4457 59814 4469 59866
rect 4521 59814 7477 59866
rect 7529 59814 7541 59866
rect 7593 59814 7605 59866
rect 7657 59814 7669 59866
rect 7721 59814 7733 59866
rect 7785 59814 10856 59866
rect 1104 59792 10856 59814
rect 1673 59619 1731 59625
rect 1673 59585 1685 59619
rect 1719 59616 1731 59619
rect 3602 59616 3608 59628
rect 1719 59588 3608 59616
rect 1719 59585 1731 59588
rect 1673 59579 1731 59585
rect 3602 59576 3608 59588
rect 3660 59576 3666 59628
rect 9858 59616 9864 59628
rect 9819 59588 9864 59616
rect 9858 59576 9864 59588
rect 9916 59576 9922 59628
rect 1394 59372 1400 59424
rect 1452 59412 1458 59424
rect 1489 59415 1547 59421
rect 1489 59412 1501 59415
rect 1452 59384 1501 59412
rect 1452 59372 1458 59384
rect 1489 59381 1501 59384
rect 1535 59381 1547 59415
rect 10042 59412 10048 59424
rect 10003 59384 10048 59412
rect 1489 59375 1547 59381
rect 10042 59372 10048 59384
rect 10100 59372 10106 59424
rect 1104 59322 10856 59344
rect 1104 59270 2582 59322
rect 2634 59270 2646 59322
rect 2698 59270 2710 59322
rect 2762 59270 2774 59322
rect 2826 59270 2838 59322
rect 2890 59270 5845 59322
rect 5897 59270 5909 59322
rect 5961 59270 5973 59322
rect 6025 59270 6037 59322
rect 6089 59270 6101 59322
rect 6153 59270 9109 59322
rect 9161 59270 9173 59322
rect 9225 59270 9237 59322
rect 9289 59270 9301 59322
rect 9353 59270 9365 59322
rect 9417 59270 10856 59322
rect 1104 59248 10856 59270
rect 1762 59100 1768 59152
rect 1820 59140 1826 59152
rect 2130 59140 2136 59152
rect 1820 59112 2136 59140
rect 1820 59100 1826 59112
rect 2130 59100 2136 59112
rect 2188 59100 2194 59152
rect 1673 59007 1731 59013
rect 1673 58973 1685 59007
rect 1719 59004 1731 59007
rect 1762 59004 1768 59016
rect 1719 58976 1768 59004
rect 1719 58973 1731 58976
rect 1673 58967 1731 58973
rect 1762 58964 1768 58976
rect 1820 58964 1826 59016
rect 1486 58868 1492 58880
rect 1447 58840 1492 58868
rect 1486 58828 1492 58840
rect 1544 58828 1550 58880
rect 1104 58778 10856 58800
rect 1104 58726 4213 58778
rect 4265 58726 4277 58778
rect 4329 58726 4341 58778
rect 4393 58726 4405 58778
rect 4457 58726 4469 58778
rect 4521 58726 7477 58778
rect 7529 58726 7541 58778
rect 7593 58726 7605 58778
rect 7657 58726 7669 58778
rect 7721 58726 7733 58778
rect 7785 58726 10856 58778
rect 1104 58704 10856 58726
rect 1673 58531 1731 58537
rect 1673 58497 1685 58531
rect 1719 58528 1731 58531
rect 1946 58528 1952 58540
rect 1719 58500 1952 58528
rect 1719 58497 1731 58500
rect 1673 58491 1731 58497
rect 1946 58488 1952 58500
rect 2004 58488 2010 58540
rect 9861 58531 9919 58537
rect 9861 58497 9873 58531
rect 9907 58528 9919 58531
rect 11517 58531 11575 58537
rect 11517 58528 11529 58531
rect 9907 58500 11529 58528
rect 9907 58497 9919 58500
rect 9861 58491 9919 58497
rect 11517 58497 11529 58500
rect 11563 58497 11575 58531
rect 11517 58491 11575 58497
rect 10042 58392 10048 58404
rect 10003 58364 10048 58392
rect 10042 58352 10048 58364
rect 10100 58352 10106 58404
rect 1394 58284 1400 58336
rect 1452 58324 1458 58336
rect 1489 58327 1547 58333
rect 1489 58324 1501 58327
rect 1452 58296 1501 58324
rect 1452 58284 1458 58296
rect 1489 58293 1501 58296
rect 1535 58293 1547 58327
rect 1489 58287 1547 58293
rect 1104 58234 10856 58256
rect 1104 58182 2582 58234
rect 2634 58182 2646 58234
rect 2698 58182 2710 58234
rect 2762 58182 2774 58234
rect 2826 58182 2838 58234
rect 2890 58182 5845 58234
rect 5897 58182 5909 58234
rect 5961 58182 5973 58234
rect 6025 58182 6037 58234
rect 6089 58182 6101 58234
rect 6153 58182 9109 58234
rect 9161 58182 9173 58234
rect 9225 58182 9237 58234
rect 9289 58182 9301 58234
rect 9353 58182 9365 58234
rect 9417 58182 10856 58234
rect 1104 58160 10856 58182
rect 1302 58012 1308 58064
rect 1360 58052 1366 58064
rect 2222 58052 2228 58064
rect 1360 58024 2228 58052
rect 1360 58012 1366 58024
rect 2222 58012 2228 58024
rect 2280 58012 2286 58064
rect 2148 57956 2544 57984
rect 1397 57919 1455 57925
rect 1397 57885 1409 57919
rect 1443 57885 1455 57919
rect 1397 57879 1455 57885
rect 1412 57780 1440 57879
rect 1486 57876 1492 57928
rect 1544 57916 1550 57928
rect 1673 57919 1731 57925
rect 1673 57916 1685 57919
rect 1544 57888 1685 57916
rect 1544 57876 1550 57888
rect 1673 57885 1685 57888
rect 1719 57885 1731 57919
rect 1673 57879 1731 57885
rect 1765 57919 1823 57925
rect 1765 57885 1777 57919
rect 1811 57916 1823 57919
rect 2148 57916 2176 57956
rect 1811 57888 2176 57916
rect 1811 57885 1823 57888
rect 1765 57879 1823 57885
rect 2222 57876 2228 57928
rect 2280 57916 2286 57928
rect 2409 57919 2467 57925
rect 2409 57916 2421 57919
rect 2280 57888 2421 57916
rect 2280 57876 2286 57888
rect 2409 57885 2421 57888
rect 2455 57885 2467 57919
rect 2516 57916 2544 57956
rect 2590 57916 2596 57928
rect 2516 57888 2596 57916
rect 2409 57879 2467 57885
rect 2590 57876 2596 57888
rect 2648 57876 2654 57928
rect 9861 57919 9919 57925
rect 9861 57885 9873 57919
rect 9907 57916 9919 57919
rect 11149 57919 11207 57925
rect 11149 57916 11161 57919
rect 9907 57888 11161 57916
rect 9907 57885 9919 57888
rect 9861 57879 9919 57885
rect 11149 57885 11161 57888
rect 11195 57885 11207 57919
rect 11149 57879 11207 57885
rect 1581 57851 1639 57857
rect 1581 57817 1593 57851
rect 1627 57817 1639 57851
rect 8570 57848 8576 57860
rect 1581 57811 1639 57817
rect 1872 57820 8576 57848
rect 1486 57780 1492 57792
rect 1412 57752 1492 57780
rect 1486 57740 1492 57752
rect 1544 57740 1550 57792
rect 1596 57780 1624 57811
rect 1872 57780 1900 57820
rect 8570 57808 8576 57820
rect 8628 57808 8634 57860
rect 1596 57752 1900 57780
rect 1946 57740 1952 57792
rect 2004 57780 2010 57792
rect 2593 57783 2651 57789
rect 2004 57752 2049 57780
rect 2004 57740 2010 57752
rect 2593 57749 2605 57783
rect 2639 57780 2651 57783
rect 2774 57780 2780 57792
rect 2639 57752 2780 57780
rect 2639 57749 2651 57752
rect 2593 57743 2651 57749
rect 2774 57740 2780 57752
rect 2832 57740 2838 57792
rect 10042 57780 10048 57792
rect 10003 57752 10048 57780
rect 10042 57740 10048 57752
rect 10100 57740 10106 57792
rect 1104 57690 10856 57712
rect 1104 57638 4213 57690
rect 4265 57638 4277 57690
rect 4329 57638 4341 57690
rect 4393 57638 4405 57690
rect 4457 57638 4469 57690
rect 4521 57638 7477 57690
rect 7529 57638 7541 57690
rect 7593 57638 7605 57690
rect 7657 57638 7669 57690
rect 7721 57638 7733 57690
rect 7785 57638 10856 57690
rect 1104 57616 10856 57638
rect 1946 57536 1952 57588
rect 2004 57576 2010 57588
rect 11057 57579 11115 57585
rect 11057 57576 11069 57579
rect 2004 57548 11069 57576
rect 2004 57536 2010 57548
rect 11057 57545 11069 57548
rect 11103 57545 11115 57579
rect 11057 57539 11115 57545
rect 1670 57508 1676 57520
rect 1631 57480 1676 57508
rect 1670 57468 1676 57480
rect 1728 57468 1734 57520
rect 3142 57468 3148 57520
rect 3200 57508 3206 57520
rect 3326 57508 3332 57520
rect 3200 57480 3332 57508
rect 3200 57468 3206 57480
rect 3326 57468 3332 57480
rect 3384 57468 3390 57520
rect 1397 57443 1455 57449
rect 1397 57409 1409 57443
rect 1443 57440 1455 57443
rect 1486 57440 1492 57452
rect 1443 57412 1492 57440
rect 1443 57409 1455 57412
rect 1397 57403 1455 57409
rect 1486 57400 1492 57412
rect 1544 57400 1550 57452
rect 1581 57443 1639 57449
rect 1581 57409 1593 57443
rect 1627 57409 1639 57443
rect 1581 57403 1639 57409
rect 1765 57443 1823 57449
rect 1765 57409 1777 57443
rect 1811 57440 1823 57443
rect 1946 57440 1952 57452
rect 1811 57412 1952 57440
rect 1811 57409 1823 57412
rect 1765 57403 1823 57409
rect 1596 57372 1624 57403
rect 1946 57400 1952 57412
rect 2004 57440 2010 57452
rect 2590 57440 2596 57452
rect 2004 57412 2596 57440
rect 2004 57400 2010 57412
rect 2590 57400 2596 57412
rect 2648 57400 2654 57452
rect 2685 57443 2743 57449
rect 2685 57409 2697 57443
rect 2731 57440 2743 57443
rect 3510 57440 3516 57452
rect 2731 57412 3516 57440
rect 2731 57409 2743 57412
rect 2685 57403 2743 57409
rect 3510 57400 3516 57412
rect 3568 57400 3574 57452
rect 9861 57443 9919 57449
rect 9861 57409 9873 57443
rect 9907 57440 9919 57443
rect 11333 57443 11391 57449
rect 11333 57440 11345 57443
rect 9907 57412 11345 57440
rect 9907 57409 9919 57412
rect 9861 57403 9919 57409
rect 11333 57409 11345 57412
rect 11379 57409 11391 57443
rect 11333 57403 11391 57409
rect 7374 57372 7380 57384
rect 1596 57344 7380 57372
rect 7374 57332 7380 57344
rect 7432 57332 7438 57384
rect 1949 57307 2007 57313
rect 1949 57273 1961 57307
rect 1995 57304 2007 57307
rect 9858 57304 9864 57316
rect 1995 57276 9864 57304
rect 1995 57273 2007 57276
rect 1949 57267 2007 57273
rect 9858 57264 9864 57276
rect 9916 57264 9922 57316
rect 2501 57239 2559 57245
rect 2501 57205 2513 57239
rect 2547 57236 2559 57239
rect 2958 57236 2964 57248
rect 2547 57208 2964 57236
rect 2547 57205 2559 57208
rect 2501 57199 2559 57205
rect 2958 57196 2964 57208
rect 3016 57196 3022 57248
rect 10042 57236 10048 57248
rect 10003 57208 10048 57236
rect 10042 57196 10048 57208
rect 10100 57196 10106 57248
rect 1104 57146 10856 57168
rect 1104 57094 2582 57146
rect 2634 57094 2646 57146
rect 2698 57094 2710 57146
rect 2762 57094 2774 57146
rect 2826 57094 2838 57146
rect 2890 57094 5845 57146
rect 5897 57094 5909 57146
rect 5961 57094 5973 57146
rect 6025 57094 6037 57146
rect 6089 57094 6101 57146
rect 6153 57094 9109 57146
rect 9161 57094 9173 57146
rect 9225 57094 9237 57146
rect 9289 57094 9301 57146
rect 9353 57094 9365 57146
rect 9417 57094 10856 57146
rect 1104 57072 10856 57094
rect 2777 57035 2835 57041
rect 2777 57001 2789 57035
rect 2823 57032 2835 57035
rect 3053 57035 3111 57041
rect 3053 57032 3065 57035
rect 2823 57004 3065 57032
rect 2823 57001 2835 57004
rect 2777 56995 2835 57001
rect 3053 57001 3065 57004
rect 3099 57032 3111 57035
rect 3234 57032 3240 57044
rect 3099 57004 3240 57032
rect 3099 57001 3111 57004
rect 3053 56995 3111 57001
rect 3234 56992 3240 57004
rect 3292 57032 3298 57044
rect 3878 57032 3884 57044
rect 3292 57004 3884 57032
rect 3292 56992 3298 57004
rect 3878 56992 3884 57004
rect 3936 56992 3942 57044
rect 1949 56967 2007 56973
rect 1949 56933 1961 56967
rect 1995 56964 2007 56967
rect 9766 56964 9772 56976
rect 1995 56936 9772 56964
rect 1995 56933 2007 56936
rect 1949 56927 2007 56933
rect 9766 56924 9772 56936
rect 9824 56924 9830 56976
rect 7282 56896 7288 56908
rect 1596 56868 7288 56896
rect 1394 56828 1400 56840
rect 1355 56800 1400 56828
rect 1394 56788 1400 56800
rect 1452 56788 1458 56840
rect 1596 56837 1624 56868
rect 7282 56856 7288 56868
rect 7340 56856 7346 56908
rect 1581 56831 1639 56837
rect 1581 56797 1593 56831
rect 1627 56797 1639 56831
rect 1581 56791 1639 56797
rect 1765 56831 1823 56837
rect 1765 56797 1777 56831
rect 1811 56828 1823 56831
rect 1946 56828 1952 56840
rect 1811 56800 1952 56828
rect 1811 56797 1823 56800
rect 1765 56791 1823 56797
rect 1946 56788 1952 56800
rect 2004 56828 2010 56840
rect 2682 56828 2688 56840
rect 2004 56800 2688 56828
rect 2004 56788 2010 56800
rect 2682 56788 2688 56800
rect 2740 56788 2746 56840
rect 3789 56831 3847 56837
rect 3789 56797 3801 56831
rect 3835 56828 3847 56831
rect 3878 56828 3884 56840
rect 3835 56800 3884 56828
rect 3835 56797 3847 56800
rect 3789 56791 3847 56797
rect 3878 56788 3884 56800
rect 3936 56788 3942 56840
rect 1673 56763 1731 56769
rect 1673 56729 1685 56763
rect 1719 56760 1731 56763
rect 2038 56760 2044 56772
rect 1719 56732 2044 56760
rect 1719 56729 1731 56732
rect 1673 56723 1731 56729
rect 2038 56720 2044 56732
rect 2096 56720 2102 56772
rect 2961 56763 3019 56769
rect 2961 56729 2973 56763
rect 3007 56760 3019 56763
rect 3142 56760 3148 56772
rect 3007 56732 3148 56760
rect 3007 56729 3019 56732
rect 2961 56723 3019 56729
rect 3142 56720 3148 56732
rect 3200 56720 3206 56772
rect 1854 56692 1860 56704
rect 1044 56664 1860 56692
rect 1044 56488 1072 56664
rect 1854 56652 1860 56664
rect 1912 56652 1918 56704
rect 1946 56652 1952 56704
rect 2004 56692 2010 56704
rect 2222 56692 2228 56704
rect 2004 56664 2228 56692
rect 2004 56652 2010 56664
rect 2222 56652 2228 56664
rect 2280 56652 2286 56704
rect 2777 56695 2835 56701
rect 2777 56661 2789 56695
rect 2823 56692 2835 56695
rect 2866 56692 2872 56704
rect 2823 56664 2872 56692
rect 2823 56661 2835 56664
rect 2777 56655 2835 56661
rect 2866 56652 2872 56664
rect 2924 56652 2930 56704
rect 3970 56692 3976 56704
rect 3931 56664 3976 56692
rect 3970 56652 3976 56664
rect 4028 56652 4034 56704
rect 1104 56602 10856 56624
rect 1104 56550 4213 56602
rect 4265 56550 4277 56602
rect 4329 56550 4341 56602
rect 4393 56550 4405 56602
rect 4457 56550 4469 56602
rect 4521 56550 7477 56602
rect 7529 56550 7541 56602
rect 7593 56550 7605 56602
rect 7657 56550 7669 56602
rect 7721 56550 7733 56602
rect 7785 56550 10856 56602
rect 1104 56528 10856 56550
rect 1044 56460 1532 56488
rect 1394 56352 1400 56364
rect 1355 56324 1400 56352
rect 1394 56312 1400 56324
rect 1452 56312 1458 56364
rect 1504 56352 1532 56460
rect 1670 56448 1676 56500
rect 1728 56488 1734 56500
rect 2590 56488 2596 56500
rect 1728 56460 2596 56488
rect 1728 56448 1734 56460
rect 2590 56448 2596 56460
rect 2648 56448 2654 56500
rect 3602 56448 3608 56500
rect 3660 56488 3666 56500
rect 3973 56491 4031 56497
rect 3660 56460 3740 56488
rect 3660 56448 3666 56460
rect 1581 56423 1639 56429
rect 1581 56389 1593 56423
rect 1627 56420 1639 56423
rect 3712 56420 3740 56460
rect 3973 56457 3985 56491
rect 4019 56488 4031 56491
rect 4062 56488 4068 56500
rect 4019 56460 4068 56488
rect 4019 56457 4031 56460
rect 3973 56451 4031 56457
rect 4062 56448 4068 56460
rect 4120 56448 4126 56500
rect 11241 56491 11299 56497
rect 11241 56457 11253 56491
rect 11287 56457 11299 56491
rect 11241 56451 11299 56457
rect 1627 56392 3004 56420
rect 3712 56392 4016 56420
rect 1627 56389 1639 56392
rect 1581 56383 1639 56389
rect 1673 56355 1731 56361
rect 1673 56352 1685 56355
rect 1504 56324 1685 56352
rect 1673 56321 1685 56324
rect 1719 56321 1731 56355
rect 1673 56315 1731 56321
rect 1765 56355 1823 56361
rect 1765 56321 1777 56355
rect 1811 56352 1823 56355
rect 2682 56352 2688 56364
rect 1811 56324 2688 56352
rect 1811 56321 1823 56324
rect 1765 56315 1823 56321
rect 1872 56160 1900 56324
rect 2682 56312 2688 56324
rect 2740 56352 2746 56364
rect 2777 56355 2835 56361
rect 2777 56352 2789 56355
rect 2740 56324 2789 56352
rect 2740 56312 2746 56324
rect 2777 56321 2789 56324
rect 2823 56321 2835 56355
rect 2777 56315 2835 56321
rect 2501 56287 2559 56293
rect 2501 56253 2513 56287
rect 2547 56284 2559 56287
rect 2866 56284 2872 56296
rect 2547 56256 2872 56284
rect 2547 56253 2559 56256
rect 2501 56247 2559 56253
rect 2866 56244 2872 56256
rect 2924 56244 2930 56296
rect 2976 56284 3004 56392
rect 3050 56312 3056 56364
rect 3108 56352 3114 56364
rect 3602 56352 3608 56364
rect 3108 56324 3608 56352
rect 3108 56312 3114 56324
rect 3602 56312 3608 56324
rect 3660 56352 3666 56364
rect 3789 56355 3847 56361
rect 3789 56352 3801 56355
rect 3660 56324 3801 56352
rect 3660 56312 3666 56324
rect 3789 56321 3801 56324
rect 3835 56321 3847 56355
rect 3789 56315 3847 56321
rect 3988 56296 4016 56392
rect 5810 56380 5816 56432
rect 5868 56420 5874 56432
rect 11256 56420 11284 56451
rect 5868 56392 11284 56420
rect 5868 56380 5874 56392
rect 9861 56355 9919 56361
rect 9861 56321 9873 56355
rect 9907 56352 9919 56355
rect 11241 56355 11299 56361
rect 11241 56352 11253 56355
rect 9907 56324 11253 56352
rect 9907 56321 9919 56324
rect 9861 56315 9919 56321
rect 11241 56321 11253 56324
rect 11287 56321 11299 56355
rect 11241 56315 11299 56321
rect 2976 56256 3924 56284
rect 1949 56219 2007 56225
rect 1949 56185 1961 56219
rect 1995 56216 2007 56219
rect 3050 56216 3056 56228
rect 1995 56188 3056 56216
rect 1995 56185 2007 56188
rect 1949 56179 2007 56185
rect 3050 56176 3056 56188
rect 3108 56176 3114 56228
rect 3896 56216 3924 56256
rect 3970 56244 3976 56296
rect 4028 56244 4034 56296
rect 8662 56216 8668 56228
rect 3896 56188 8668 56216
rect 8662 56176 8668 56188
rect 8720 56176 8726 56228
rect 1854 56108 1860 56160
rect 1912 56108 1918 56160
rect 10042 56148 10048 56160
rect 10003 56120 10048 56148
rect 10042 56108 10048 56120
rect 10100 56108 10106 56160
rect 1104 56058 10856 56080
rect 1104 56006 2582 56058
rect 2634 56006 2646 56058
rect 2698 56006 2710 56058
rect 2762 56006 2774 56058
rect 2826 56006 2838 56058
rect 2890 56006 5845 56058
rect 5897 56006 5909 56058
rect 5961 56006 5973 56058
rect 6025 56006 6037 56058
rect 6089 56006 6101 56058
rect 6153 56006 9109 56058
rect 9161 56006 9173 56058
rect 9225 56006 9237 56058
rect 9289 56006 9301 56058
rect 9353 56006 9365 56058
rect 9417 56006 10856 56058
rect 1104 55984 10856 56006
rect 1394 55768 1400 55820
rect 1452 55808 1458 55820
rect 2225 55811 2283 55817
rect 2225 55808 2237 55811
rect 1452 55780 2237 55808
rect 1452 55768 1458 55780
rect 2225 55777 2237 55780
rect 2271 55777 2283 55811
rect 2225 55771 2283 55777
rect 4062 55768 4068 55820
rect 4120 55768 4126 55820
rect 1949 55743 2007 55749
rect 1949 55709 1961 55743
rect 1995 55709 2007 55743
rect 1949 55703 2007 55709
rect 1964 55672 1992 55703
rect 2314 55700 2320 55752
rect 2372 55740 2378 55752
rect 3789 55743 3847 55749
rect 3789 55740 3801 55743
rect 2372 55712 3801 55740
rect 2372 55700 2378 55712
rect 3789 55709 3801 55712
rect 3835 55709 3847 55743
rect 3789 55703 3847 55709
rect 3050 55672 3056 55684
rect 1964 55644 3056 55672
rect 3050 55632 3056 55644
rect 3108 55672 3114 55684
rect 4080 55672 4108 55768
rect 9861 55743 9919 55749
rect 9861 55709 9873 55743
rect 9907 55740 9919 55743
rect 11057 55743 11115 55749
rect 11057 55740 11069 55743
rect 9907 55712 11069 55740
rect 9907 55709 9919 55712
rect 9861 55703 9919 55709
rect 11057 55709 11069 55712
rect 11103 55709 11115 55743
rect 11057 55703 11115 55709
rect 3108 55644 4108 55672
rect 3108 55632 3114 55644
rect 3970 55604 3976 55616
rect 3931 55576 3976 55604
rect 3970 55564 3976 55576
rect 4028 55564 4034 55616
rect 10042 55604 10048 55616
rect 10003 55576 10048 55604
rect 10042 55564 10048 55576
rect 10100 55564 10106 55616
rect 1104 55514 10856 55536
rect 1104 55462 4213 55514
rect 4265 55462 4277 55514
rect 4329 55462 4341 55514
rect 4393 55462 4405 55514
rect 4457 55462 4469 55514
rect 4521 55462 7477 55514
rect 7529 55462 7541 55514
rect 7593 55462 7605 55514
rect 7657 55462 7669 55514
rect 7721 55462 7733 55514
rect 7785 55462 10856 55514
rect 1104 55440 10856 55462
rect 1949 55403 2007 55409
rect 1949 55369 1961 55403
rect 1995 55400 2007 55403
rect 1995 55372 2636 55400
rect 1995 55369 2007 55372
rect 1949 55363 2007 55369
rect 1581 55335 1639 55341
rect 1581 55301 1593 55335
rect 1627 55332 1639 55335
rect 2608 55332 2636 55372
rect 2682 55360 2688 55412
rect 2740 55400 2746 55412
rect 2958 55400 2964 55412
rect 2740 55372 2964 55400
rect 2740 55360 2746 55372
rect 2958 55360 2964 55372
rect 3016 55360 3022 55412
rect 11425 55335 11483 55341
rect 11425 55332 11437 55335
rect 1627 55304 2544 55332
rect 2608 55304 11437 55332
rect 1627 55301 1639 55304
rect 1581 55295 1639 55301
rect 1394 55264 1400 55276
rect 1355 55236 1400 55264
rect 1394 55224 1400 55236
rect 1452 55224 1458 55276
rect 1670 55264 1676 55276
rect 1631 55236 1676 55264
rect 1670 55224 1676 55236
rect 1728 55224 1734 55276
rect 1765 55267 1823 55273
rect 1765 55233 1777 55267
rect 1811 55264 1823 55267
rect 1854 55264 1860 55276
rect 1811 55236 1860 55264
rect 1811 55233 1823 55236
rect 1765 55227 1823 55233
rect 1854 55224 1860 55236
rect 1912 55224 1918 55276
rect 2038 55224 2044 55276
rect 2096 55264 2102 55276
rect 2409 55267 2467 55273
rect 2409 55264 2421 55267
rect 2096 55236 2421 55264
rect 2096 55224 2102 55236
rect 2409 55233 2421 55236
rect 2455 55233 2467 55267
rect 2516 55264 2544 55304
rect 11425 55301 11437 55304
rect 11471 55301 11483 55335
rect 11425 55295 11483 55301
rect 8754 55264 8760 55276
rect 2516 55236 8760 55264
rect 2409 55227 2467 55233
rect 8754 55224 8760 55236
rect 8812 55224 8818 55276
rect 1578 55156 1584 55208
rect 1636 55156 1642 55208
rect 4706 55156 4712 55208
rect 4764 55196 4770 55208
rect 5534 55196 5540 55208
rect 4764 55168 5540 55196
rect 4764 55156 4770 55168
rect 5534 55156 5540 55168
rect 5592 55156 5598 55208
rect 1394 55088 1400 55140
rect 1452 55128 1458 55140
rect 1596 55128 1624 55156
rect 1452 55100 1624 55128
rect 2593 55131 2651 55137
rect 1452 55088 1458 55100
rect 2593 55097 2605 55131
rect 2639 55128 2651 55131
rect 2682 55128 2688 55140
rect 2639 55100 2688 55128
rect 2639 55097 2651 55100
rect 2593 55091 2651 55097
rect 2682 55088 2688 55100
rect 2740 55088 2746 55140
rect 1104 54970 10856 54992
rect 1104 54918 2582 54970
rect 2634 54918 2646 54970
rect 2698 54918 2710 54970
rect 2762 54918 2774 54970
rect 2826 54918 2838 54970
rect 2890 54918 5845 54970
rect 5897 54918 5909 54970
rect 5961 54918 5973 54970
rect 6025 54918 6037 54970
rect 6089 54918 6101 54970
rect 6153 54918 9109 54970
rect 9161 54918 9173 54970
rect 9225 54918 9237 54970
rect 9289 54918 9301 54970
rect 9353 54918 9365 54970
rect 9417 54918 10856 54970
rect 1104 54896 10856 54918
rect 1394 54612 1400 54664
rect 1452 54652 1458 54664
rect 1673 54655 1731 54661
rect 1673 54652 1685 54655
rect 1452 54624 1685 54652
rect 1452 54612 1458 54624
rect 1673 54621 1685 54624
rect 1719 54621 1731 54655
rect 10134 54652 10140 54664
rect 10095 54624 10140 54652
rect 1673 54615 1731 54621
rect 10134 54612 10140 54624
rect 10192 54612 10198 54664
rect 1486 54516 1492 54528
rect 1447 54488 1492 54516
rect 1486 54476 1492 54488
rect 1544 54476 1550 54528
rect 9950 54516 9956 54528
rect 9911 54488 9956 54516
rect 9950 54476 9956 54488
rect 10008 54476 10014 54528
rect 1104 54426 10856 54448
rect 1104 54374 4213 54426
rect 4265 54374 4277 54426
rect 4329 54374 4341 54426
rect 4393 54374 4405 54426
rect 4457 54374 4469 54426
rect 4521 54374 7477 54426
rect 7529 54374 7541 54426
rect 7593 54374 7605 54426
rect 7657 54374 7669 54426
rect 7721 54374 7733 54426
rect 7785 54374 10856 54426
rect 1104 54352 10856 54374
rect 3142 54204 3148 54256
rect 3200 54244 3206 54256
rect 3789 54247 3847 54253
rect 3789 54244 3801 54247
rect 3200 54216 3801 54244
rect 3200 54204 3206 54216
rect 3789 54213 3801 54216
rect 3835 54213 3847 54247
rect 3789 54207 3847 54213
rect 845 54179 903 54185
rect 845 54145 857 54179
rect 891 54176 903 54179
rect 1673 54179 1731 54185
rect 1673 54176 1685 54179
rect 891 54148 1685 54176
rect 891 54145 903 54148
rect 845 54139 903 54145
rect 1673 54145 1685 54148
rect 1719 54145 1731 54179
rect 1673 54139 1731 54145
rect 2501 54179 2559 54185
rect 2501 54145 2513 54179
rect 2547 54176 2559 54179
rect 3234 54176 3240 54188
rect 2547 54148 3240 54176
rect 2547 54145 2559 54148
rect 2501 54139 2559 54145
rect 3234 54136 3240 54148
rect 3292 54136 3298 54188
rect 3970 54176 3976 54188
rect 3931 54148 3976 54176
rect 3970 54136 3976 54148
rect 4028 54136 4034 54188
rect 10134 54176 10140 54188
rect 10095 54148 10140 54176
rect 10134 54136 10140 54148
rect 10192 54136 10198 54188
rect 2777 54111 2835 54117
rect 2777 54077 2789 54111
rect 2823 54108 2835 54111
rect 2958 54108 2964 54120
rect 2823 54080 2964 54108
rect 2823 54077 2835 54080
rect 2777 54071 2835 54077
rect 2958 54068 2964 54080
rect 3016 54068 3022 54120
rect 3142 54068 3148 54120
rect 3200 54108 3206 54120
rect 3510 54108 3516 54120
rect 3200 54080 3516 54108
rect 3200 54068 3206 54080
rect 3510 54068 3516 54080
rect 3568 54068 3574 54120
rect 1486 53972 1492 53984
rect 1447 53944 1492 53972
rect 1486 53932 1492 53944
rect 1544 53932 1550 53984
rect 9858 53932 9864 53984
rect 9916 53972 9922 53984
rect 9953 53975 10011 53981
rect 9953 53972 9965 53975
rect 9916 53944 9965 53972
rect 9916 53932 9922 53944
rect 9953 53941 9965 53944
rect 9999 53941 10011 53975
rect 9953 53935 10011 53941
rect 1104 53882 10856 53904
rect 1104 53830 2582 53882
rect 2634 53830 2646 53882
rect 2698 53830 2710 53882
rect 2762 53830 2774 53882
rect 2826 53830 2838 53882
rect 2890 53830 5845 53882
rect 5897 53830 5909 53882
rect 5961 53830 5973 53882
rect 6025 53830 6037 53882
rect 6089 53830 6101 53882
rect 6153 53830 9109 53882
rect 9161 53830 9173 53882
rect 9225 53830 9237 53882
rect 9289 53830 9301 53882
rect 9353 53830 9365 53882
rect 9417 53830 10856 53882
rect 1104 53808 10856 53830
rect 2041 53635 2099 53641
rect 2041 53601 2053 53635
rect 2087 53632 2099 53635
rect 3050 53632 3056 53644
rect 2087 53604 3056 53632
rect 2087 53601 2099 53604
rect 2041 53595 2099 53601
rect 3050 53592 3056 53604
rect 3108 53592 3114 53644
rect 2222 53524 2228 53576
rect 2280 53564 2286 53576
rect 2317 53567 2375 53573
rect 2317 53564 2329 53567
rect 2280 53536 2329 53564
rect 2280 53524 2286 53536
rect 2317 53533 2329 53536
rect 2363 53533 2375 53567
rect 2317 53527 2375 53533
rect 6733 53567 6791 53573
rect 6733 53533 6745 53567
rect 6779 53564 6791 53567
rect 9950 53564 9956 53576
rect 6779 53536 9956 53564
rect 6779 53533 6791 53536
rect 6733 53527 6791 53533
rect 9950 53524 9956 53536
rect 10008 53524 10014 53576
rect 10134 53564 10140 53576
rect 10095 53536 10140 53564
rect 10134 53524 10140 53536
rect 10192 53524 10198 53576
rect 3050 53388 3056 53440
rect 3108 53428 3114 53440
rect 6549 53431 6607 53437
rect 6549 53428 6561 53431
rect 3108 53400 6561 53428
rect 3108 53388 3114 53400
rect 6549 53397 6561 53400
rect 6595 53397 6607 53431
rect 9950 53428 9956 53440
rect 9911 53400 9956 53428
rect 6549 53391 6607 53397
rect 9950 53388 9956 53400
rect 10008 53388 10014 53440
rect 1104 53338 10856 53360
rect 1104 53286 4213 53338
rect 4265 53286 4277 53338
rect 4329 53286 4341 53338
rect 4393 53286 4405 53338
rect 4457 53286 4469 53338
rect 4521 53286 7477 53338
rect 7529 53286 7541 53338
rect 7593 53286 7605 53338
rect 7657 53286 7669 53338
rect 7721 53286 7733 53338
rect 7785 53286 10856 53338
rect 1104 53264 10856 53286
rect 1486 53184 1492 53236
rect 1544 53224 1550 53236
rect 2317 53227 2375 53233
rect 2317 53224 2329 53227
rect 1544 53196 2329 53224
rect 1544 53184 1550 53196
rect 2317 53193 2329 53196
rect 2363 53193 2375 53227
rect 2317 53187 2375 53193
rect 2961 53227 3019 53233
rect 2961 53193 2973 53227
rect 3007 53224 3019 53227
rect 3786 53224 3792 53236
rect 3007 53196 3792 53224
rect 3007 53193 3019 53196
rect 2961 53187 3019 53193
rect 3786 53184 3792 53196
rect 3844 53184 3850 53236
rect 842 53116 848 53168
rect 900 53156 906 53168
rect 900 53128 3096 53156
rect 900 53116 906 53128
rect 3068 53100 3096 53128
rect 1673 53091 1731 53097
rect 1673 53057 1685 53091
rect 1719 53057 1731 53091
rect 1673 53051 1731 53057
rect 1688 53020 1716 53051
rect 1946 53048 1952 53100
rect 2004 53088 2010 53100
rect 2133 53091 2191 53097
rect 2133 53088 2145 53091
rect 2004 53060 2145 53088
rect 2004 53048 2010 53060
rect 2133 53057 2145 53060
rect 2179 53057 2191 53091
rect 2133 53051 2191 53057
rect 2774 53048 2780 53100
rect 2832 53088 2838 53100
rect 2869 53091 2927 53097
rect 2869 53088 2881 53091
rect 2832 53060 2881 53088
rect 2832 53048 2838 53060
rect 2869 53057 2881 53060
rect 2915 53057 2927 53091
rect 3050 53088 3056 53100
rect 3011 53060 3056 53088
rect 2869 53051 2927 53057
rect 3050 53048 3056 53060
rect 3108 53048 3114 53100
rect 7193 53091 7251 53097
rect 7193 53057 7205 53091
rect 7239 53088 7251 53091
rect 9858 53088 9864 53100
rect 7239 53060 9864 53088
rect 7239 53057 7251 53060
rect 7193 53051 7251 53057
rect 9858 53048 9864 53060
rect 9916 53048 9922 53100
rect 3510 53020 3516 53032
rect 1688 52992 3516 53020
rect 3510 52980 3516 52992
rect 3568 52980 3574 53032
rect 198 52912 204 52964
rect 256 52952 262 52964
rect 256 52924 1624 52952
rect 256 52912 262 52924
rect 1486 52884 1492 52896
rect 1447 52856 1492 52884
rect 1486 52844 1492 52856
rect 1544 52844 1550 52896
rect 1596 52884 1624 52924
rect 3234 52884 3240 52896
rect 1596 52856 3240 52884
rect 3234 52844 3240 52856
rect 3292 52884 3298 52896
rect 7101 52887 7159 52893
rect 7101 52884 7113 52887
rect 3292 52856 7113 52884
rect 3292 52844 3298 52856
rect 7101 52853 7113 52856
rect 7147 52853 7159 52887
rect 7101 52847 7159 52853
rect 1104 52794 10856 52816
rect 1104 52742 2582 52794
rect 2634 52742 2646 52794
rect 2698 52742 2710 52794
rect 2762 52742 2774 52794
rect 2826 52742 2838 52794
rect 2890 52742 5845 52794
rect 5897 52742 5909 52794
rect 5961 52742 5973 52794
rect 6025 52742 6037 52794
rect 6089 52742 6101 52794
rect 6153 52742 9109 52794
rect 9161 52742 9173 52794
rect 9225 52742 9237 52794
rect 9289 52742 9301 52794
rect 9353 52742 9365 52794
rect 9417 52742 10856 52794
rect 1104 52720 10856 52742
rect 1302 52640 1308 52692
rect 1360 52680 1366 52692
rect 1670 52680 1676 52692
rect 1360 52652 1676 52680
rect 1360 52640 1366 52652
rect 1670 52640 1676 52652
rect 1728 52640 1734 52692
rect 2406 52680 2412 52692
rect 2367 52652 2412 52680
rect 2406 52640 2412 52652
rect 2464 52640 2470 52692
rect 3053 52683 3111 52689
rect 3053 52649 3065 52683
rect 3099 52680 3111 52683
rect 3694 52680 3700 52692
rect 3099 52652 3700 52680
rect 3099 52649 3111 52652
rect 3053 52643 3111 52649
rect 3694 52640 3700 52652
rect 3752 52640 3758 52692
rect 750 52572 756 52624
rect 808 52612 814 52624
rect 9033 52615 9091 52621
rect 9033 52612 9045 52615
rect 808 52584 9045 52612
rect 808 52572 814 52584
rect 2516 52544 2544 52584
rect 9033 52581 9045 52584
rect 9079 52581 9091 52615
rect 9033 52575 9091 52581
rect 3142 52544 3148 52556
rect 2516 52516 2636 52544
rect 2608 52485 2636 52516
rect 3068 52516 3148 52544
rect 3068 52485 3096 52516
rect 3142 52504 3148 52516
rect 3200 52504 3206 52556
rect 1673 52479 1731 52485
rect 1673 52445 1685 52479
rect 1719 52476 1731 52479
rect 2409 52479 2467 52485
rect 1719 52448 2360 52476
rect 1719 52445 1731 52448
rect 1673 52439 1731 52445
rect 1486 52340 1492 52352
rect 1447 52312 1492 52340
rect 1486 52300 1492 52312
rect 1544 52300 1550 52352
rect 2332 52340 2360 52448
rect 2409 52445 2421 52479
rect 2455 52445 2467 52479
rect 2409 52439 2467 52445
rect 2587 52479 2645 52485
rect 2587 52445 2599 52479
rect 2633 52445 2645 52479
rect 2587 52439 2645 52445
rect 3053 52479 3111 52485
rect 3053 52445 3065 52479
rect 3099 52445 3111 52479
rect 3234 52476 3240 52488
rect 3195 52448 3240 52476
rect 3053 52439 3111 52445
rect 2424 52408 2452 52439
rect 3068 52408 3096 52439
rect 3234 52436 3240 52448
rect 3292 52436 3298 52488
rect 9125 52479 9183 52485
rect 9125 52445 9137 52479
rect 9171 52476 9183 52479
rect 9950 52476 9956 52488
rect 9171 52448 9956 52476
rect 9171 52445 9183 52448
rect 9125 52439 9183 52445
rect 9950 52436 9956 52448
rect 10008 52436 10014 52488
rect 10134 52476 10140 52488
rect 10095 52448 10140 52476
rect 10134 52436 10140 52448
rect 10192 52436 10198 52488
rect 5442 52408 5448 52420
rect 2424 52380 5448 52408
rect 5442 52368 5448 52380
rect 5500 52368 5506 52420
rect 3142 52340 3148 52352
rect 2332 52312 3148 52340
rect 3142 52300 3148 52312
rect 3200 52300 3206 52352
rect 3602 52300 3608 52352
rect 3660 52340 3666 52352
rect 4062 52340 4068 52352
rect 3660 52312 4068 52340
rect 3660 52300 3666 52312
rect 4062 52300 4068 52312
rect 4120 52300 4126 52352
rect 9490 52300 9496 52352
rect 9548 52340 9554 52352
rect 9953 52343 10011 52349
rect 9953 52340 9965 52343
rect 9548 52312 9965 52340
rect 9548 52300 9554 52312
rect 9953 52309 9965 52312
rect 9999 52309 10011 52343
rect 9953 52303 10011 52309
rect 1104 52250 10856 52272
rect 1104 52198 4213 52250
rect 4265 52198 4277 52250
rect 4329 52198 4341 52250
rect 4393 52198 4405 52250
rect 4457 52198 4469 52250
rect 4521 52198 7477 52250
rect 7529 52198 7541 52250
rect 7593 52198 7605 52250
rect 7657 52198 7669 52250
rect 7721 52198 7733 52250
rect 7785 52198 10856 52250
rect 1104 52176 10856 52198
rect 2130 52136 2136 52148
rect 1504 52108 2136 52136
rect 1397 52003 1455 52009
rect 1397 51969 1409 52003
rect 1443 51969 1455 52003
rect 1504 52000 1532 52108
rect 2130 52096 2136 52108
rect 2188 52096 2194 52148
rect 3237 52139 3295 52145
rect 3237 52105 3249 52139
rect 3283 52136 3295 52139
rect 3418 52136 3424 52148
rect 3283 52108 3424 52136
rect 3283 52105 3295 52108
rect 3237 52099 3295 52105
rect 3418 52096 3424 52108
rect 3476 52096 3482 52148
rect 1581 52071 1639 52077
rect 1581 52037 1593 52071
rect 1627 52068 1639 52071
rect 8018 52068 8024 52080
rect 1627 52040 8024 52068
rect 1627 52037 1639 52040
rect 1581 52031 1639 52037
rect 8018 52028 8024 52040
rect 8076 52028 8082 52080
rect 1673 52003 1731 52009
rect 1673 52000 1685 52003
rect 1504 51972 1685 52000
rect 1397 51963 1455 51969
rect 1673 51969 1685 51972
rect 1719 51969 1731 52003
rect 1673 51963 1731 51969
rect 1765 52003 1823 52009
rect 1765 51969 1777 52003
rect 1811 52000 1823 52003
rect 2130 52000 2136 52012
rect 1811 51972 2136 52000
rect 1811 51969 1823 51972
rect 1765 51963 1823 51969
rect 1412 51796 1440 51963
rect 2130 51960 2136 51972
rect 2188 51960 2194 52012
rect 2409 52003 2467 52009
rect 2409 51969 2421 52003
rect 2455 52000 2467 52003
rect 2498 52000 2504 52012
rect 2455 51972 2504 52000
rect 2455 51969 2467 51972
rect 2409 51963 2467 51969
rect 2498 51960 2504 51972
rect 2556 51960 2562 52012
rect 3145 52003 3203 52009
rect 3145 51969 3157 52003
rect 3191 51969 3203 52003
rect 3145 51963 3203 51969
rect 3329 52003 3387 52009
rect 3329 51969 3341 52003
rect 3375 52000 3387 52003
rect 4062 52000 4068 52012
rect 3375 51972 4068 52000
rect 3375 51969 3387 51972
rect 3329 51963 3387 51969
rect 3160 51932 3188 51963
rect 4062 51960 4068 51972
rect 4120 51960 4126 52012
rect 10134 52000 10140 52012
rect 10095 51972 10140 52000
rect 10134 51960 10140 51972
rect 10192 51960 10198 52012
rect 3418 51932 3424 51944
rect 3160 51904 3424 51932
rect 3418 51892 3424 51904
rect 3476 51892 3482 51944
rect 1949 51867 2007 51873
rect 1949 51833 1961 51867
rect 1995 51864 2007 51867
rect 2593 51867 2651 51873
rect 1995 51836 2360 51864
rect 1995 51833 2007 51836
rect 1949 51827 2007 51833
rect 2222 51796 2228 51808
rect 1412 51768 2228 51796
rect 2222 51756 2228 51768
rect 2280 51756 2286 51808
rect 2332 51796 2360 51836
rect 2593 51833 2605 51867
rect 2639 51864 2651 51867
rect 2774 51864 2780 51876
rect 2639 51836 2780 51864
rect 2639 51833 2651 51836
rect 2593 51827 2651 51833
rect 2774 51824 2780 51836
rect 2832 51824 2838 51876
rect 11057 51867 11115 51873
rect 11057 51864 11069 51867
rect 3068 51836 11069 51864
rect 3068 51796 3096 51836
rect 11057 51833 11069 51836
rect 11103 51833 11115 51867
rect 11057 51827 11115 51833
rect 9950 51796 9956 51808
rect 2332 51768 3096 51796
rect 9911 51768 9956 51796
rect 9950 51756 9956 51768
rect 10008 51756 10014 51808
rect 1104 51706 10856 51728
rect 1104 51654 2582 51706
rect 2634 51654 2646 51706
rect 2698 51654 2710 51706
rect 2762 51654 2774 51706
rect 2826 51654 2838 51706
rect 2890 51654 5845 51706
rect 5897 51654 5909 51706
rect 5961 51654 5973 51706
rect 6025 51654 6037 51706
rect 6089 51654 6101 51706
rect 6153 51654 9109 51706
rect 9161 51654 9173 51706
rect 9225 51654 9237 51706
rect 9289 51654 9301 51706
rect 9353 51654 9365 51706
rect 9417 51654 10856 51706
rect 1104 51632 10856 51654
rect 2406 51592 2412 51604
rect 1596 51564 2412 51592
rect 937 51459 995 51465
rect 937 51425 949 51459
rect 983 51456 995 51459
rect 983 51428 1532 51456
rect 983 51425 995 51428
rect 937 51419 995 51425
rect 1397 51391 1455 51397
rect 1397 51357 1409 51391
rect 1443 51357 1455 51391
rect 1397 51351 1455 51357
rect 1412 51252 1440 51351
rect 1504 51264 1532 51428
rect 1596 51397 1624 51564
rect 2406 51552 2412 51564
rect 2464 51552 2470 51604
rect 2961 51595 3019 51601
rect 2961 51561 2973 51595
rect 3007 51592 3019 51595
rect 11149 51595 11207 51601
rect 11149 51592 11161 51595
rect 3007 51564 11161 51592
rect 3007 51561 3019 51564
rect 2961 51555 3019 51561
rect 11149 51561 11161 51564
rect 11195 51561 11207 51595
rect 11149 51555 11207 51561
rect 1949 51527 2007 51533
rect 1949 51493 1961 51527
rect 1995 51524 2007 51527
rect 2590 51524 2596 51536
rect 1995 51496 2596 51524
rect 1995 51493 2007 51496
rect 1949 51487 2007 51493
rect 2590 51484 2596 51496
rect 2648 51484 2654 51536
rect 2130 51456 2136 51468
rect 1826 51428 2136 51456
rect 1581 51391 1639 51397
rect 1581 51357 1593 51391
rect 1627 51357 1639 51391
rect 1581 51351 1639 51357
rect 1670 51348 1676 51400
rect 1728 51388 1734 51400
rect 1826 51397 1854 51428
rect 2130 51416 2136 51428
rect 2188 51456 2194 51468
rect 2314 51456 2320 51468
rect 2188 51428 2320 51456
rect 2188 51416 2194 51428
rect 2314 51416 2320 51428
rect 2372 51456 2378 51468
rect 2372 51428 2820 51456
rect 2372 51416 2378 51428
rect 1811 51391 1869 51397
rect 1728 51360 1773 51388
rect 1728 51348 1734 51360
rect 1811 51357 1823 51391
rect 1857 51357 1869 51391
rect 1811 51351 1869 51357
rect 2222 51348 2228 51400
rect 2280 51388 2286 51400
rect 2406 51388 2412 51400
rect 2280 51360 2412 51388
rect 2280 51348 2286 51360
rect 2406 51348 2412 51360
rect 2464 51348 2470 51400
rect 2792 51397 2820 51428
rect 5810 51416 5816 51468
rect 5868 51456 5874 51468
rect 11241 51459 11299 51465
rect 11241 51456 11253 51459
rect 5868 51428 11253 51456
rect 5868 51416 5874 51428
rect 11241 51425 11253 51428
rect 11287 51425 11299 51459
rect 11241 51419 11299 51425
rect 2777 51391 2835 51397
rect 2777 51357 2789 51391
rect 2823 51388 2835 51391
rect 2958 51388 2964 51400
rect 2823 51360 2964 51388
rect 2823 51357 2835 51360
rect 2777 51351 2835 51357
rect 2958 51348 2964 51360
rect 3016 51348 3022 51400
rect 3234 51348 3240 51400
rect 3292 51348 3298 51400
rect 4341 51391 4399 51397
rect 4341 51357 4353 51391
rect 4387 51388 4399 51391
rect 9490 51388 9496 51400
rect 4387 51360 9496 51388
rect 4387 51357 4399 51360
rect 4341 51351 4399 51357
rect 9490 51348 9496 51360
rect 9548 51348 9554 51400
rect 2593 51323 2651 51329
rect 2593 51289 2605 51323
rect 2639 51289 2651 51323
rect 2593 51283 2651 51289
rect 2685 51323 2743 51329
rect 2685 51289 2697 51323
rect 2731 51320 2743 51323
rect 3252 51320 3280 51348
rect 2731 51292 3280 51320
rect 2731 51289 2743 51292
rect 2685 51283 2743 51289
rect 1044 51224 1440 51252
rect 1044 51048 1072 51224
rect 1486 51212 1492 51264
rect 1544 51212 1550 51264
rect 1578 51212 1584 51264
rect 1636 51252 1642 51264
rect 2130 51252 2136 51264
rect 1636 51224 2136 51252
rect 1636 51212 1642 51224
rect 2130 51212 2136 51224
rect 2188 51212 2194 51264
rect 2608 51252 2636 51283
rect 3234 51252 3240 51264
rect 2608 51224 3240 51252
rect 3234 51212 3240 51224
rect 3292 51212 3298 51264
rect 4157 51255 4215 51261
rect 4157 51221 4169 51255
rect 4203 51252 4215 51255
rect 4890 51252 4896 51264
rect 4203 51224 4896 51252
rect 4203 51221 4215 51224
rect 4157 51215 4215 51221
rect 4890 51212 4896 51224
rect 4948 51212 4954 51264
rect 1104 51162 10856 51184
rect 1104 51110 4213 51162
rect 4265 51110 4277 51162
rect 4329 51110 4341 51162
rect 4393 51110 4405 51162
rect 4457 51110 4469 51162
rect 4521 51110 7477 51162
rect 7529 51110 7541 51162
rect 7593 51110 7605 51162
rect 7657 51110 7669 51162
rect 7721 51110 7733 51162
rect 7785 51110 10856 51162
rect 1104 51088 10856 51110
rect 2406 51048 2412 51060
rect 1044 51020 2412 51048
rect 1412 50924 1440 51020
rect 2406 51008 2412 51020
rect 2464 51008 2470 51060
rect 3237 51051 3295 51057
rect 3237 51017 3249 51051
rect 3283 51048 3295 51051
rect 3602 51048 3608 51060
rect 3283 51020 3608 51048
rect 3283 51017 3295 51020
rect 3237 51011 3295 51017
rect 3602 51008 3608 51020
rect 3660 51008 3666 51060
rect 9950 51048 9956 51060
rect 4080 51020 9956 51048
rect 1670 50980 1676 50992
rect 1631 50952 1676 50980
rect 1670 50940 1676 50952
rect 1728 50940 1734 50992
rect 2314 50980 2320 50992
rect 1780 50952 2320 50980
rect 1394 50912 1400 50924
rect 1307 50884 1400 50912
rect 1394 50872 1400 50884
rect 1452 50872 1458 50924
rect 1780 50921 1808 50952
rect 2314 50940 2320 50952
rect 2372 50940 2378 50992
rect 1581 50915 1639 50921
rect 1581 50881 1593 50915
rect 1627 50881 1639 50915
rect 1581 50875 1639 50881
rect 1765 50915 1823 50921
rect 1765 50881 1777 50915
rect 1811 50881 1823 50915
rect 2406 50912 2412 50924
rect 2367 50884 2412 50912
rect 1765 50875 1823 50881
rect 1596 50844 1624 50875
rect 2406 50872 2412 50884
rect 2464 50872 2470 50924
rect 3145 50915 3203 50921
rect 3145 50881 3157 50915
rect 3191 50881 3203 50915
rect 3145 50875 3203 50881
rect 3329 50915 3387 50921
rect 3329 50881 3341 50915
rect 3375 50912 3387 50915
rect 3528 50912 3648 50916
rect 3712 50912 3924 50916
rect 3970 50912 3976 50924
rect 3375 50888 3976 50912
rect 3375 50884 3556 50888
rect 3620 50884 3740 50888
rect 3896 50884 3976 50888
rect 3375 50881 3387 50884
rect 3329 50875 3387 50881
rect 3050 50844 3056 50856
rect 1596 50816 3056 50844
rect 3050 50804 3056 50816
rect 3108 50804 3114 50856
rect 3160 50844 3188 50875
rect 3970 50872 3976 50884
rect 4028 50872 4034 50924
rect 4080 50921 4108 51020
rect 9950 51008 9956 51020
rect 10008 51008 10014 51060
rect 4065 50915 4123 50921
rect 4065 50881 4077 50915
rect 4111 50881 4123 50915
rect 4065 50875 4123 50881
rect 4709 50915 4767 50921
rect 4709 50881 4721 50915
rect 4755 50881 4767 50915
rect 4890 50912 4896 50924
rect 4851 50884 4896 50912
rect 4709 50875 4767 50881
rect 4724 50844 4752 50875
rect 4890 50872 4896 50884
rect 4948 50872 4954 50924
rect 10134 50912 10140 50924
rect 10095 50884 10140 50912
rect 10134 50872 10140 50884
rect 10192 50872 10198 50924
rect 3160 50816 3372 50844
rect 3344 50788 3372 50816
rect 3804 50816 4752 50844
rect 2593 50779 2651 50785
rect 2593 50745 2605 50779
rect 2639 50776 2651 50779
rect 2774 50776 2780 50788
rect 2639 50748 2780 50776
rect 2639 50745 2651 50748
rect 2593 50739 2651 50745
rect 2774 50736 2780 50748
rect 2832 50736 2838 50788
rect 3326 50736 3332 50788
rect 3384 50776 3390 50788
rect 3804 50776 3832 50816
rect 11333 50779 11391 50785
rect 11333 50776 11345 50779
rect 3384 50748 3832 50776
rect 3896 50748 11345 50776
rect 3384 50736 3390 50748
rect 1949 50711 2007 50717
rect 1949 50677 1961 50711
rect 1995 50708 2007 50711
rect 3896 50708 3924 50748
rect 11333 50745 11345 50748
rect 11379 50745 11391 50779
rect 11333 50739 11391 50745
rect 4062 50708 4068 50720
rect 1995 50680 3924 50708
rect 4023 50680 4068 50708
rect 1995 50677 2007 50680
rect 1949 50671 2007 50677
rect 4062 50668 4068 50680
rect 4120 50668 4126 50720
rect 4154 50668 4160 50720
rect 4212 50708 4218 50720
rect 4709 50711 4767 50717
rect 4709 50708 4721 50711
rect 4212 50680 4721 50708
rect 4212 50668 4218 50680
rect 4709 50677 4721 50680
rect 4755 50677 4767 50711
rect 9950 50708 9956 50720
rect 9911 50680 9956 50708
rect 4709 50671 4767 50677
rect 9950 50668 9956 50680
rect 10008 50668 10014 50720
rect 1104 50618 10856 50640
rect 1104 50566 2582 50618
rect 2634 50566 2646 50618
rect 2698 50566 2710 50618
rect 2762 50566 2774 50618
rect 2826 50566 2838 50618
rect 2890 50566 5845 50618
rect 5897 50566 5909 50618
rect 5961 50566 5973 50618
rect 6025 50566 6037 50618
rect 6089 50566 6101 50618
rect 6153 50566 9109 50618
rect 9161 50566 9173 50618
rect 9225 50566 9237 50618
rect 9289 50566 9301 50618
rect 9353 50566 9365 50618
rect 9417 50566 10856 50618
rect 1104 50544 10856 50566
rect 3050 50464 3056 50516
rect 3108 50504 3114 50516
rect 8110 50504 8116 50516
rect 3108 50476 8116 50504
rect 3108 50464 3114 50476
rect 8110 50464 8116 50476
rect 8168 50464 8174 50516
rect 1949 50439 2007 50445
rect 1949 50405 1961 50439
rect 1995 50436 2007 50439
rect 11517 50439 11575 50445
rect 11517 50436 11529 50439
rect 1995 50408 11529 50436
rect 1995 50405 2007 50408
rect 1949 50399 2007 50405
rect 11517 50405 11529 50408
rect 11563 50405 11575 50439
rect 11517 50399 11575 50405
rect 3418 50328 3424 50380
rect 3476 50368 3482 50380
rect 4154 50368 4160 50380
rect 3476 50340 4160 50368
rect 3476 50328 3482 50340
rect 4154 50328 4160 50340
rect 4212 50328 4218 50380
rect 1394 50300 1400 50312
rect 1355 50272 1400 50300
rect 1394 50260 1400 50272
rect 1452 50260 1458 50312
rect 1486 50260 1492 50312
rect 1544 50300 1550 50312
rect 1673 50303 1731 50309
rect 1673 50300 1685 50303
rect 1544 50272 1685 50300
rect 1544 50260 1550 50272
rect 1673 50269 1685 50272
rect 1719 50269 1731 50303
rect 1673 50263 1731 50269
rect 1765 50303 1823 50309
rect 1765 50269 1777 50303
rect 1811 50300 1823 50303
rect 2314 50300 2320 50312
rect 1811 50272 2320 50300
rect 1811 50269 1823 50272
rect 1765 50263 1823 50269
rect 2314 50260 2320 50272
rect 2372 50260 2378 50312
rect 2685 50303 2743 50309
rect 2685 50269 2697 50303
rect 2731 50300 2743 50303
rect 3050 50300 3056 50312
rect 2731 50272 3056 50300
rect 2731 50269 2743 50272
rect 2685 50263 2743 50269
rect 3050 50260 3056 50272
rect 3108 50260 3114 50312
rect 4249 50303 4307 50309
rect 4249 50269 4261 50303
rect 4295 50300 4307 50303
rect 9950 50300 9956 50312
rect 4295 50272 9956 50300
rect 4295 50269 4307 50272
rect 4249 50263 4307 50269
rect 9950 50260 9956 50272
rect 10008 50260 10014 50312
rect 10134 50300 10140 50312
rect 10095 50272 10140 50300
rect 10134 50260 10140 50272
rect 10192 50260 10198 50312
rect 1581 50235 1639 50241
rect 1581 50201 1593 50235
rect 1627 50201 1639 50235
rect 3418 50232 3424 50244
rect 1581 50195 1639 50201
rect 1872 50204 3424 50232
rect 1596 50164 1624 50195
rect 1872 50164 1900 50204
rect 3418 50192 3424 50204
rect 3476 50192 3482 50244
rect 2498 50164 2504 50176
rect 1596 50136 1900 50164
rect 2459 50136 2504 50164
rect 2498 50124 2504 50136
rect 2556 50124 2562 50176
rect 3970 50124 3976 50176
rect 4028 50164 4034 50176
rect 4065 50167 4123 50173
rect 4065 50164 4077 50167
rect 4028 50136 4077 50164
rect 4028 50124 4034 50136
rect 4065 50133 4077 50136
rect 4111 50164 4123 50167
rect 6270 50164 6276 50176
rect 4111 50136 6276 50164
rect 4111 50133 4123 50136
rect 4065 50127 4123 50133
rect 6270 50124 6276 50136
rect 6328 50124 6334 50176
rect 9950 50164 9956 50176
rect 9911 50136 9956 50164
rect 9950 50124 9956 50136
rect 10008 50124 10014 50176
rect 1104 50074 10856 50096
rect 1104 50022 4213 50074
rect 4265 50022 4277 50074
rect 4329 50022 4341 50074
rect 4393 50022 4405 50074
rect 4457 50022 4469 50074
rect 4521 50022 7477 50074
rect 7529 50022 7541 50074
rect 7593 50022 7605 50074
rect 7657 50022 7669 50074
rect 7721 50022 7733 50074
rect 7785 50022 10856 50074
rect 1104 50000 10856 50022
rect 1762 49920 1768 49972
rect 1820 49960 1826 49972
rect 2409 49963 2467 49969
rect 2409 49960 2421 49963
rect 1820 49932 2421 49960
rect 1820 49920 1826 49932
rect 2409 49929 2421 49932
rect 2455 49929 2467 49963
rect 4065 49963 4123 49969
rect 4065 49960 4077 49963
rect 2409 49923 2467 49929
rect 2746 49932 4077 49960
rect 1673 49827 1731 49833
rect 1673 49793 1685 49827
rect 1719 49824 1731 49827
rect 1762 49824 1768 49836
rect 1719 49796 1768 49824
rect 1719 49793 1731 49796
rect 1673 49787 1731 49793
rect 1762 49784 1768 49796
rect 1820 49784 1826 49836
rect 2317 49827 2375 49833
rect 2317 49793 2329 49827
rect 2363 49793 2375 49827
rect 2317 49787 2375 49793
rect 2501 49827 2559 49833
rect 2501 49793 2513 49827
rect 2547 49824 2559 49827
rect 2746 49824 2774 49932
rect 4065 49929 4077 49932
rect 4111 49960 4123 49963
rect 4706 49960 4712 49972
rect 4111 49932 4712 49960
rect 4111 49929 4123 49932
rect 4065 49923 4123 49929
rect 4706 49920 4712 49932
rect 4764 49920 4770 49972
rect 2547 49796 2774 49824
rect 3421 49827 3479 49833
rect 2547 49793 2559 49796
rect 2501 49787 2559 49793
rect 3421 49793 3433 49827
rect 3467 49824 3479 49827
rect 3510 49824 3516 49836
rect 3467 49796 3516 49824
rect 3467 49793 3479 49796
rect 3421 49787 3479 49793
rect 1486 49688 1492 49700
rect 1447 49660 1492 49688
rect 1486 49648 1492 49660
rect 1544 49648 1550 49700
rect 2332 49688 2360 49787
rect 3510 49784 3516 49796
rect 3568 49824 3574 49836
rect 3970 49824 3976 49836
rect 3568 49796 3976 49824
rect 3568 49784 3574 49796
rect 3970 49784 3976 49796
rect 4028 49784 4034 49836
rect 4249 49827 4307 49833
rect 4249 49793 4261 49827
rect 4295 49824 4307 49827
rect 9950 49824 9956 49836
rect 4295 49796 9956 49824
rect 4295 49793 4307 49796
rect 4249 49787 4307 49793
rect 9950 49784 9956 49796
rect 10008 49784 10014 49836
rect 10137 49827 10195 49833
rect 10137 49793 10149 49827
rect 10183 49793 10195 49827
rect 10137 49787 10195 49793
rect 4062 49716 4068 49768
rect 4120 49756 4126 49768
rect 4982 49756 4988 49768
rect 4120 49728 4988 49756
rect 4120 49716 4126 49728
rect 4982 49716 4988 49728
rect 5040 49716 5046 49768
rect 10152 49700 10180 49787
rect 3326 49688 3332 49700
rect 2332 49660 3332 49688
rect 3326 49648 3332 49660
rect 3384 49648 3390 49700
rect 5442 49688 5448 49700
rect 3436 49660 5448 49688
rect 3237 49623 3295 49629
rect 3237 49589 3249 49623
rect 3283 49620 3295 49623
rect 3436 49620 3464 49660
rect 5442 49648 5448 49660
rect 5500 49648 5506 49700
rect 10134 49648 10140 49700
rect 10192 49648 10198 49700
rect 3283 49592 3464 49620
rect 3283 49589 3295 49592
rect 3237 49583 3295 49589
rect 4246 49580 4252 49632
rect 4304 49620 4310 49632
rect 9953 49623 10011 49629
rect 9953 49620 9965 49623
rect 4304 49592 9965 49620
rect 4304 49580 4310 49592
rect 9953 49589 9965 49592
rect 9999 49589 10011 49623
rect 9953 49583 10011 49589
rect 1104 49530 10856 49552
rect 1104 49478 2582 49530
rect 2634 49478 2646 49530
rect 2698 49478 2710 49530
rect 2762 49478 2774 49530
rect 2826 49478 2838 49530
rect 2890 49478 5845 49530
rect 5897 49478 5909 49530
rect 5961 49478 5973 49530
rect 6025 49478 6037 49530
rect 6089 49478 6101 49530
rect 6153 49478 9109 49530
rect 9161 49478 9173 49530
rect 9225 49478 9237 49530
rect 9289 49478 9301 49530
rect 9353 49478 9365 49530
rect 9417 49478 10856 49530
rect 1104 49456 10856 49478
rect 1854 49376 1860 49428
rect 1912 49416 1918 49428
rect 2317 49419 2375 49425
rect 2317 49416 2329 49419
rect 1912 49388 2329 49416
rect 1912 49376 1918 49388
rect 2317 49385 2329 49388
rect 2363 49385 2375 49419
rect 2317 49379 2375 49385
rect 658 49240 664 49292
rect 716 49280 722 49292
rect 3973 49283 4031 49289
rect 3973 49280 3985 49283
rect 716 49252 3985 49280
rect 716 49240 722 49252
rect 1673 49215 1731 49221
rect 1673 49181 1685 49215
rect 1719 49212 1731 49215
rect 1854 49212 1860 49224
rect 1719 49184 1860 49212
rect 1719 49181 1731 49184
rect 1673 49175 1731 49181
rect 1854 49172 1860 49184
rect 1912 49172 1918 49224
rect 2516 49221 2544 49252
rect 3973 49249 3985 49252
rect 4019 49249 4031 49283
rect 3973 49243 4031 49249
rect 2317 49215 2375 49221
rect 2317 49181 2329 49215
rect 2363 49181 2375 49215
rect 2317 49175 2375 49181
rect 2501 49215 2559 49221
rect 2501 49181 2513 49215
rect 2547 49212 2559 49215
rect 4246 49212 4252 49224
rect 2547 49184 2581 49212
rect 4207 49184 4252 49212
rect 2547 49181 2559 49184
rect 2501 49175 2559 49181
rect 2332 49144 2360 49175
rect 4246 49172 4252 49184
rect 4304 49172 4310 49224
rect 3326 49144 3332 49156
rect 2332 49116 3332 49144
rect 3326 49104 3332 49116
rect 3384 49104 3390 49156
rect 1486 49076 1492 49088
rect 1447 49048 1492 49076
rect 1486 49036 1492 49048
rect 1544 49036 1550 49088
rect 1104 48986 10856 49008
rect 1104 48934 4213 48986
rect 4265 48934 4277 48986
rect 4329 48934 4341 48986
rect 4393 48934 4405 48986
rect 4457 48934 4469 48986
rect 4521 48934 7477 48986
rect 7529 48934 7541 48986
rect 7593 48934 7605 48986
rect 7657 48934 7669 48986
rect 7721 48934 7733 48986
rect 7785 48934 10856 48986
rect 1104 48912 10856 48934
rect 3786 48872 3792 48884
rect 3747 48844 3792 48872
rect 3786 48832 3792 48844
rect 3844 48832 3850 48884
rect 1673 48739 1731 48745
rect 1673 48705 1685 48739
rect 1719 48736 1731 48739
rect 3510 48736 3516 48748
rect 1719 48708 3516 48736
rect 1719 48705 1731 48708
rect 1673 48699 1731 48705
rect 3510 48696 3516 48708
rect 3568 48696 3574 48748
rect 3973 48739 4031 48745
rect 3973 48705 3985 48739
rect 4019 48705 4031 48739
rect 10134 48736 10140 48748
rect 10095 48708 10140 48736
rect 3973 48699 4031 48705
rect 566 48628 572 48680
rect 624 48668 630 48680
rect 3988 48668 4016 48699
rect 10134 48696 10140 48708
rect 10192 48696 10198 48748
rect 624 48640 4016 48668
rect 624 48628 630 48640
rect 1486 48600 1492 48612
rect 1447 48572 1492 48600
rect 1486 48560 1492 48572
rect 1544 48560 1550 48612
rect 845 48535 903 48541
rect 845 48501 857 48535
rect 891 48532 903 48535
rect 3786 48532 3792 48544
rect 891 48504 3792 48532
rect 891 48501 903 48504
rect 845 48495 903 48501
rect 3786 48492 3792 48504
rect 3844 48492 3850 48544
rect 9950 48532 9956 48544
rect 9911 48504 9956 48532
rect 9950 48492 9956 48504
rect 10008 48492 10014 48544
rect 1104 48442 10856 48464
rect 1104 48390 2582 48442
rect 2634 48390 2646 48442
rect 2698 48390 2710 48442
rect 2762 48390 2774 48442
rect 2826 48390 2838 48442
rect 2890 48390 5845 48442
rect 5897 48390 5909 48442
rect 5961 48390 5973 48442
rect 6025 48390 6037 48442
rect 6089 48390 6101 48442
rect 6153 48390 9109 48442
rect 9161 48390 9173 48442
rect 9225 48390 9237 48442
rect 9289 48390 9301 48442
rect 9353 48390 9365 48442
rect 9417 48390 10856 48442
rect 1104 48368 10856 48390
rect 1673 48127 1731 48133
rect 1673 48093 1685 48127
rect 1719 48124 1731 48127
rect 2314 48124 2320 48136
rect 1719 48096 2320 48124
rect 1719 48093 1731 48096
rect 1673 48087 1731 48093
rect 2314 48084 2320 48096
rect 2372 48084 2378 48136
rect 10134 48124 10140 48136
rect 10095 48096 10140 48124
rect 10134 48084 10140 48096
rect 10192 48084 10198 48136
rect 1486 47988 1492 48000
rect 1447 47960 1492 47988
rect 1486 47948 1492 47960
rect 1544 47948 1550 48000
rect 9858 47948 9864 48000
rect 9916 47988 9922 48000
rect 9953 47991 10011 47997
rect 9953 47988 9965 47991
rect 9916 47960 9965 47988
rect 9916 47948 9922 47960
rect 9953 47957 9965 47960
rect 9999 47957 10011 47991
rect 9953 47951 10011 47957
rect 1104 47898 10856 47920
rect 1104 47846 4213 47898
rect 4265 47846 4277 47898
rect 4329 47846 4341 47898
rect 4393 47846 4405 47898
rect 4457 47846 4469 47898
rect 4521 47846 7477 47898
rect 7529 47846 7541 47898
rect 7593 47846 7605 47898
rect 7657 47846 7669 47898
rect 7721 47846 7733 47898
rect 7785 47846 10856 47898
rect 1104 47824 10856 47846
rect 750 47608 756 47660
rect 808 47608 814 47660
rect 1670 47648 1676 47660
rect 1631 47620 1676 47648
rect 1670 47608 1676 47620
rect 1728 47608 1734 47660
rect 3326 47648 3332 47660
rect 3287 47620 3332 47648
rect 3326 47608 3332 47620
rect 3384 47608 3390 47660
rect 4341 47651 4399 47657
rect 4341 47617 4353 47651
rect 4387 47648 4399 47651
rect 9950 47648 9956 47660
rect 4387 47620 9956 47648
rect 4387 47617 4399 47620
rect 4341 47611 4399 47617
rect 9950 47608 9956 47620
rect 10008 47608 10014 47660
rect 768 47444 796 47608
rect 3602 47580 3608 47592
rect 3563 47552 3608 47580
rect 3602 47540 3608 47552
rect 3660 47540 3666 47592
rect 1486 47512 1492 47524
rect 1447 47484 1492 47512
rect 1486 47472 1492 47484
rect 1544 47472 1550 47524
rect 842 47444 848 47456
rect 768 47416 848 47444
rect 842 47404 848 47416
rect 900 47404 906 47456
rect 4154 47444 4160 47456
rect 4115 47416 4160 47444
rect 4154 47404 4160 47416
rect 4212 47404 4218 47456
rect 1104 47354 10856 47376
rect 1104 47302 2582 47354
rect 2634 47302 2646 47354
rect 2698 47302 2710 47354
rect 2762 47302 2774 47354
rect 2826 47302 2838 47354
rect 2890 47302 5845 47354
rect 5897 47302 5909 47354
rect 5961 47302 5973 47354
rect 6025 47302 6037 47354
rect 6089 47302 6101 47354
rect 6153 47302 9109 47354
rect 9161 47302 9173 47354
rect 9225 47302 9237 47354
rect 9289 47302 9301 47354
rect 9353 47302 9365 47354
rect 9417 47302 10856 47354
rect 1104 47280 10856 47302
rect 1486 47172 1492 47184
rect 1447 47144 1492 47172
rect 1486 47132 1492 47144
rect 1544 47132 1550 47184
rect 1673 47039 1731 47045
rect 1673 47005 1685 47039
rect 1719 47036 1731 47039
rect 3326 47036 3332 47048
rect 1719 47008 3332 47036
rect 1719 47005 1731 47008
rect 1673 46999 1731 47005
rect 3326 46996 3332 47008
rect 3384 46996 3390 47048
rect 10134 47036 10140 47048
rect 10095 47008 10140 47036
rect 10134 46996 10140 47008
rect 10192 46996 10198 47048
rect 4062 46860 4068 46912
rect 4120 46900 4126 46912
rect 9953 46903 10011 46909
rect 9953 46900 9965 46903
rect 4120 46872 9965 46900
rect 4120 46860 4126 46872
rect 9953 46869 9965 46872
rect 9999 46869 10011 46903
rect 9953 46863 10011 46869
rect 1104 46810 10856 46832
rect 1104 46758 4213 46810
rect 4265 46758 4277 46810
rect 4329 46758 4341 46810
rect 4393 46758 4405 46810
rect 4457 46758 4469 46810
rect 4521 46758 7477 46810
rect 7529 46758 7541 46810
rect 7593 46758 7605 46810
rect 7657 46758 7669 46810
rect 7721 46758 7733 46810
rect 7785 46758 10856 46810
rect 1104 46736 10856 46758
rect 2130 46656 2136 46708
rect 2188 46696 2194 46708
rect 2225 46699 2283 46705
rect 2225 46696 2237 46699
rect 2188 46668 2237 46696
rect 2188 46656 2194 46668
rect 2225 46665 2237 46668
rect 2271 46665 2283 46699
rect 2225 46659 2283 46665
rect 3970 46628 3976 46640
rect 2746 46600 3976 46628
rect 1578 46520 1584 46572
rect 1636 46560 1642 46572
rect 1673 46563 1731 46569
rect 1673 46560 1685 46563
rect 1636 46532 1685 46560
rect 1636 46520 1642 46532
rect 1673 46529 1685 46532
rect 1719 46529 1731 46563
rect 2130 46560 2136 46572
rect 2091 46532 2136 46560
rect 1673 46523 1731 46529
rect 2130 46520 2136 46532
rect 2188 46520 2194 46572
rect 2317 46563 2375 46569
rect 2317 46529 2329 46563
rect 2363 46560 2375 46563
rect 2746 46560 2774 46600
rect 3970 46588 3976 46600
rect 4028 46588 4034 46640
rect 2363 46532 2774 46560
rect 3697 46563 3755 46569
rect 2363 46529 2375 46532
rect 2317 46523 2375 46529
rect 3697 46529 3709 46563
rect 3743 46560 3755 46563
rect 9858 46560 9864 46572
rect 3743 46532 9864 46560
rect 3743 46529 3755 46532
rect 3697 46523 3755 46529
rect 106 46452 112 46504
rect 164 46492 170 46504
rect 2332 46492 2360 46523
rect 9858 46520 9864 46532
rect 9916 46520 9922 46572
rect 10134 46560 10140 46572
rect 10095 46532 10140 46560
rect 10134 46520 10140 46532
rect 10192 46520 10198 46572
rect 164 46464 2360 46492
rect 164 46452 170 46464
rect 3697 46427 3755 46433
rect 3697 46393 3709 46427
rect 3743 46424 3755 46427
rect 3970 46424 3976 46436
rect 3743 46396 3976 46424
rect 3743 46393 3755 46396
rect 3697 46387 3755 46393
rect 3970 46384 3976 46396
rect 4028 46424 4034 46436
rect 7926 46424 7932 46436
rect 4028 46396 7932 46424
rect 4028 46384 4034 46396
rect 7926 46384 7932 46396
rect 7984 46384 7990 46436
rect 1486 46356 1492 46368
rect 1447 46328 1492 46356
rect 1486 46316 1492 46328
rect 1544 46316 1550 46368
rect 7098 46316 7104 46368
rect 7156 46356 7162 46368
rect 7374 46356 7380 46368
rect 7156 46328 7380 46356
rect 7156 46316 7162 46328
rect 7374 46316 7380 46328
rect 7432 46316 7438 46368
rect 9950 46356 9956 46368
rect 9911 46328 9956 46356
rect 9950 46316 9956 46328
rect 10008 46316 10014 46368
rect 1104 46266 10856 46288
rect 1104 46214 2582 46266
rect 2634 46214 2646 46266
rect 2698 46214 2710 46266
rect 2762 46214 2774 46266
rect 2826 46214 2838 46266
rect 2890 46214 5845 46266
rect 5897 46214 5909 46266
rect 5961 46214 5973 46266
rect 6025 46214 6037 46266
rect 6089 46214 6101 46266
rect 6153 46214 9109 46266
rect 9161 46214 9173 46266
rect 9225 46214 9237 46266
rect 9289 46214 9301 46266
rect 9353 46214 9365 46266
rect 9417 46214 10856 46266
rect 1104 46192 10856 46214
rect 2133 46155 2191 46161
rect 2133 46121 2145 46155
rect 2179 46152 2191 46155
rect 2222 46152 2228 46164
rect 2179 46124 2228 46152
rect 2179 46121 2191 46124
rect 2133 46115 2191 46121
rect 2222 46112 2228 46124
rect 2280 46112 2286 46164
rect 2961 46155 3019 46161
rect 2961 46121 2973 46155
rect 3007 46152 3019 46155
rect 3878 46152 3884 46164
rect 3007 46124 3884 46152
rect 3007 46121 3019 46124
rect 2961 46115 3019 46121
rect 3878 46112 3884 46124
rect 3936 46112 3942 46164
rect 3510 46044 3516 46096
rect 3568 46084 3574 46096
rect 3694 46084 3700 46096
rect 3568 46056 3700 46084
rect 3568 46044 3574 46056
rect 3694 46044 3700 46056
rect 3752 46044 3758 46096
rect 7834 46044 7840 46096
rect 7892 46084 7898 46096
rect 8110 46084 8116 46096
rect 7892 46056 8116 46084
rect 7892 46044 7898 46056
rect 8110 46044 8116 46056
rect 8168 46044 8174 46096
rect 3970 46016 3976 46028
rect 2148 45988 2452 46016
rect 2148 45960 2176 45988
rect 1673 45951 1731 45957
rect 1673 45917 1685 45951
rect 1719 45917 1731 45951
rect 2130 45948 2136 45960
rect 2091 45920 2136 45948
rect 1673 45911 1731 45917
rect 1688 45880 1716 45911
rect 2130 45908 2136 45920
rect 2188 45908 2194 45960
rect 2317 45951 2375 45957
rect 2317 45917 2329 45951
rect 2363 45917 2375 45951
rect 2317 45911 2375 45917
rect 2222 45880 2228 45892
rect 1688 45852 2228 45880
rect 2222 45840 2228 45852
rect 2280 45840 2286 45892
rect 1486 45812 1492 45824
rect 1447 45784 1492 45812
rect 1486 45772 1492 45784
rect 1544 45772 1550 45824
rect 2332 45812 2360 45911
rect 2424 45880 2452 45988
rect 2792 45988 3976 46016
rect 2792 45957 2820 45988
rect 3970 45976 3976 45988
rect 4028 45976 4034 46028
rect 2777 45951 2835 45957
rect 2777 45917 2789 45951
rect 2823 45917 2835 45951
rect 2777 45911 2835 45917
rect 2961 45951 3019 45957
rect 2961 45917 2973 45951
rect 3007 45917 3019 45951
rect 2961 45911 3019 45917
rect 2590 45880 2596 45892
rect 2424 45852 2596 45880
rect 2590 45840 2596 45852
rect 2648 45880 2654 45892
rect 2976 45880 3004 45911
rect 3050 45908 3056 45960
rect 3108 45948 3114 45960
rect 3510 45948 3516 45960
rect 3108 45920 3516 45948
rect 3108 45908 3114 45920
rect 3510 45908 3516 45920
rect 3568 45908 3574 45960
rect 4062 45948 4068 45960
rect 4023 45920 4068 45948
rect 4062 45908 4068 45920
rect 4120 45908 4126 45960
rect 10134 45948 10140 45960
rect 10095 45920 10140 45948
rect 10134 45908 10140 45920
rect 10192 45908 10198 45960
rect 3786 45880 3792 45892
rect 2648 45852 3004 45880
rect 3747 45852 3792 45880
rect 2648 45840 2654 45852
rect 3786 45840 3792 45852
rect 3844 45840 3850 45892
rect 3970 45812 3976 45824
rect 2332 45784 3976 45812
rect 3970 45772 3976 45784
rect 4028 45772 4034 45824
rect 9858 45772 9864 45824
rect 9916 45812 9922 45824
rect 9953 45815 10011 45821
rect 9953 45812 9965 45815
rect 9916 45784 9965 45812
rect 9916 45772 9922 45784
rect 9953 45781 9965 45784
rect 9999 45781 10011 45815
rect 9953 45775 10011 45781
rect 1104 45722 10856 45744
rect 1104 45670 4213 45722
rect 4265 45670 4277 45722
rect 4329 45670 4341 45722
rect 4393 45670 4405 45722
rect 4457 45670 4469 45722
rect 4521 45670 7477 45722
rect 7529 45670 7541 45722
rect 7593 45670 7605 45722
rect 7657 45670 7669 45722
rect 7721 45670 7733 45722
rect 7785 45670 10856 45722
rect 1104 45648 10856 45670
rect 845 45543 903 45549
rect 845 45509 857 45543
rect 891 45540 903 45543
rect 2498 45540 2504 45552
rect 891 45512 2504 45540
rect 891 45509 903 45512
rect 845 45503 903 45509
rect 2498 45500 2504 45512
rect 2556 45500 2562 45552
rect 1394 45432 1400 45484
rect 1452 45472 1458 45484
rect 1673 45475 1731 45481
rect 1673 45472 1685 45475
rect 1452 45444 1685 45472
rect 1452 45432 1458 45444
rect 1673 45441 1685 45444
rect 1719 45441 1731 45475
rect 1673 45435 1731 45441
rect 2590 45432 2596 45484
rect 2648 45472 2654 45484
rect 2961 45475 3019 45481
rect 2961 45472 2973 45475
rect 2648 45444 2973 45472
rect 2648 45432 2654 45444
rect 2961 45441 2973 45444
rect 3007 45441 3019 45475
rect 2961 45435 3019 45441
rect 4249 45475 4307 45481
rect 4249 45441 4261 45475
rect 4295 45472 4307 45475
rect 9950 45472 9956 45484
rect 4295 45444 9956 45472
rect 4295 45441 4307 45444
rect 4249 45435 4307 45441
rect 9950 45432 9956 45444
rect 10008 45432 10014 45484
rect 2682 45404 2688 45416
rect 2643 45376 2688 45404
rect 2682 45364 2688 45376
rect 2740 45404 2746 45416
rect 4062 45404 4068 45416
rect 2740 45376 4068 45404
rect 2740 45364 2746 45376
rect 4062 45364 4068 45376
rect 4120 45364 4126 45416
rect 1486 45268 1492 45280
rect 1447 45240 1492 45268
rect 1486 45228 1492 45240
rect 1544 45228 1550 45280
rect 3970 45228 3976 45280
rect 4028 45268 4034 45280
rect 4065 45271 4123 45277
rect 4065 45268 4077 45271
rect 4028 45240 4077 45268
rect 4028 45228 4034 45240
rect 4065 45237 4077 45240
rect 4111 45268 4123 45271
rect 6730 45268 6736 45280
rect 4111 45240 6736 45268
rect 4111 45237 4123 45240
rect 4065 45231 4123 45237
rect 6730 45228 6736 45240
rect 6788 45228 6794 45280
rect 1104 45178 10856 45200
rect 1104 45126 2582 45178
rect 2634 45126 2646 45178
rect 2698 45126 2710 45178
rect 2762 45126 2774 45178
rect 2826 45126 2838 45178
rect 2890 45126 5845 45178
rect 5897 45126 5909 45178
rect 5961 45126 5973 45178
rect 6025 45126 6037 45178
rect 6089 45126 6101 45178
rect 6153 45126 9109 45178
rect 9161 45126 9173 45178
rect 9225 45126 9237 45178
rect 9289 45126 9301 45178
rect 9353 45126 9365 45178
rect 9417 45126 10856 45178
rect 1104 45104 10856 45126
rect 2038 45024 2044 45076
rect 2096 45064 2102 45076
rect 2133 45067 2191 45073
rect 2133 45064 2145 45067
rect 2096 45036 2145 45064
rect 2096 45024 2102 45036
rect 2133 45033 2145 45036
rect 2179 45033 2191 45067
rect 2133 45027 2191 45033
rect 2777 45067 2835 45073
rect 2777 45033 2789 45067
rect 2823 45064 2835 45067
rect 2958 45064 2964 45076
rect 2823 45036 2964 45064
rect 2823 45033 2835 45036
rect 2777 45027 2835 45033
rect 2958 45024 2964 45036
rect 3016 45024 3022 45076
rect 14 44956 20 45008
rect 72 44996 78 45008
rect 72 44968 2360 44996
rect 72 44956 78 44968
rect 1673 44863 1731 44869
rect 1673 44829 1685 44863
rect 1719 44829 1731 44863
rect 2130 44860 2136 44872
rect 2091 44832 2136 44860
rect 1673 44823 1731 44829
rect 1688 44792 1716 44823
rect 2130 44820 2136 44832
rect 2188 44820 2194 44872
rect 2332 44869 2360 44968
rect 2498 44888 2504 44940
rect 2556 44928 2562 44940
rect 2556 44900 2820 44928
rect 2556 44888 2562 44900
rect 2792 44869 2820 44900
rect 2317 44863 2375 44869
rect 2317 44829 2329 44863
rect 2363 44860 2375 44863
rect 2777 44863 2835 44869
rect 2363 44832 2452 44860
rect 2363 44829 2375 44832
rect 2317 44823 2375 44829
rect 2424 44792 2452 44832
rect 2777 44829 2789 44863
rect 2823 44829 2835 44863
rect 2777 44823 2835 44829
rect 2961 44863 3019 44869
rect 2961 44829 2973 44863
rect 3007 44860 3019 44863
rect 3786 44860 3792 44872
rect 3007 44832 3792 44860
rect 3007 44829 3019 44832
rect 2961 44823 3019 44829
rect 3786 44820 3792 44832
rect 3844 44860 3850 44872
rect 4249 44863 4307 44869
rect 3844 44832 4200 44860
rect 3844 44820 3850 44832
rect 3973 44795 4031 44801
rect 3973 44792 3985 44795
rect 1688 44764 2360 44792
rect 2424 44764 3985 44792
rect 1486 44724 1492 44736
rect 1447 44696 1492 44724
rect 1486 44684 1492 44696
rect 1544 44684 1550 44736
rect 1854 44684 1860 44736
rect 1912 44724 1918 44736
rect 2130 44724 2136 44736
rect 1912 44696 2136 44724
rect 1912 44684 1918 44696
rect 2130 44684 2136 44696
rect 2188 44684 2194 44736
rect 2332 44724 2360 44764
rect 3973 44761 3985 44764
rect 4019 44761 4031 44795
rect 4172 44792 4200 44832
rect 4249 44829 4261 44863
rect 4295 44860 4307 44863
rect 9858 44860 9864 44872
rect 4295 44832 9864 44860
rect 4295 44829 4307 44832
rect 4249 44823 4307 44829
rect 9858 44820 9864 44832
rect 9916 44820 9922 44872
rect 10134 44860 10140 44872
rect 10095 44832 10140 44860
rect 10134 44820 10140 44832
rect 10192 44820 10198 44872
rect 6362 44792 6368 44804
rect 4172 44764 6368 44792
rect 3973 44755 4031 44761
rect 6362 44752 6368 44764
rect 6420 44752 6426 44804
rect 2774 44724 2780 44736
rect 2332 44696 2780 44724
rect 2774 44684 2780 44696
rect 2832 44684 2838 44736
rect 3510 44684 3516 44736
rect 3568 44724 3574 44736
rect 3786 44724 3792 44736
rect 3568 44696 3792 44724
rect 3568 44684 3574 44696
rect 3786 44684 3792 44696
rect 3844 44684 3850 44736
rect 9950 44724 9956 44736
rect 9911 44696 9956 44724
rect 9950 44684 9956 44696
rect 10008 44684 10014 44736
rect 1104 44634 10856 44656
rect 1104 44582 4213 44634
rect 4265 44582 4277 44634
rect 4329 44582 4341 44634
rect 4393 44582 4405 44634
rect 4457 44582 4469 44634
rect 4521 44582 7477 44634
rect 7529 44582 7541 44634
rect 7593 44582 7605 44634
rect 7657 44582 7669 44634
rect 7721 44582 7733 44634
rect 7785 44582 10856 44634
rect 1104 44560 10856 44582
rect 1673 44387 1731 44393
rect 1673 44353 1685 44387
rect 1719 44384 1731 44387
rect 10134 44384 10140 44396
rect 1719 44356 2084 44384
rect 10095 44356 10140 44384
rect 1719 44353 1731 44356
rect 1673 44347 1731 44353
rect 2056 44328 2084 44356
rect 10134 44344 10140 44356
rect 10192 44344 10198 44396
rect 2038 44276 2044 44328
rect 2096 44276 2102 44328
rect 1486 44180 1492 44192
rect 1447 44152 1492 44180
rect 1486 44140 1492 44152
rect 1544 44140 1550 44192
rect 9858 44140 9864 44192
rect 9916 44180 9922 44192
rect 9953 44183 10011 44189
rect 9953 44180 9965 44183
rect 9916 44152 9965 44180
rect 9916 44140 9922 44152
rect 9953 44149 9965 44152
rect 9999 44149 10011 44183
rect 9953 44143 10011 44149
rect 1104 44090 10856 44112
rect 1104 44038 2582 44090
rect 2634 44038 2646 44090
rect 2698 44038 2710 44090
rect 2762 44038 2774 44090
rect 2826 44038 2838 44090
rect 2890 44038 5845 44090
rect 5897 44038 5909 44090
rect 5961 44038 5973 44090
rect 6025 44038 6037 44090
rect 6089 44038 6101 44090
rect 6153 44038 9109 44090
rect 9161 44038 9173 44090
rect 9225 44038 9237 44090
rect 9289 44038 9301 44090
rect 9353 44038 9365 44090
rect 9417 44038 10856 44090
rect 1104 44016 10856 44038
rect 1673 43775 1731 43781
rect 1673 43741 1685 43775
rect 1719 43772 1731 43775
rect 2498 43772 2504 43784
rect 1719 43744 2504 43772
rect 1719 43741 1731 43744
rect 1673 43735 1731 43741
rect 2498 43732 2504 43744
rect 2556 43732 2562 43784
rect 10134 43772 10140 43784
rect 10095 43744 10140 43772
rect 10134 43732 10140 43744
rect 10192 43732 10198 43784
rect 1486 43636 1492 43648
rect 1447 43608 1492 43636
rect 1486 43596 1492 43608
rect 1544 43596 1550 43648
rect 9766 43596 9772 43648
rect 9824 43636 9830 43648
rect 9953 43639 10011 43645
rect 9953 43636 9965 43639
rect 9824 43608 9965 43636
rect 9824 43596 9830 43608
rect 9953 43605 9965 43608
rect 9999 43605 10011 43639
rect 9953 43599 10011 43605
rect 1104 43546 10856 43568
rect 1104 43494 4213 43546
rect 4265 43494 4277 43546
rect 4329 43494 4341 43546
rect 4393 43494 4405 43546
rect 4457 43494 4469 43546
rect 4521 43494 7477 43546
rect 7529 43494 7541 43546
rect 7593 43494 7605 43546
rect 7657 43494 7669 43546
rect 7721 43494 7733 43546
rect 7785 43494 10856 43546
rect 1104 43472 10856 43494
rect 1673 43299 1731 43305
rect 1673 43265 1685 43299
rect 1719 43296 1731 43299
rect 3326 43296 3332 43308
rect 1719 43268 3332 43296
rect 1719 43265 1731 43268
rect 1673 43259 1731 43265
rect 3326 43256 3332 43268
rect 3384 43256 3390 43308
rect 3789 43299 3847 43305
rect 3789 43265 3801 43299
rect 3835 43296 3847 43299
rect 9950 43296 9956 43308
rect 3835 43268 9956 43296
rect 3835 43265 3847 43268
rect 3789 43259 3847 43265
rect 9950 43256 9956 43268
rect 10008 43256 10014 43308
rect 1486 43092 1492 43104
rect 1447 43064 1492 43092
rect 1486 43052 1492 43064
rect 1544 43052 1550 43104
rect 3510 43052 3516 43104
rect 3568 43092 3574 43104
rect 3605 43095 3663 43101
rect 3605 43092 3617 43095
rect 3568 43064 3617 43092
rect 3568 43052 3574 43064
rect 3605 43061 3617 43064
rect 3651 43061 3663 43095
rect 3605 43055 3663 43061
rect 1104 43002 10856 43024
rect 1104 42950 2582 43002
rect 2634 42950 2646 43002
rect 2698 42950 2710 43002
rect 2762 42950 2774 43002
rect 2826 42950 2838 43002
rect 2890 42950 5845 43002
rect 5897 42950 5909 43002
rect 5961 42950 5973 43002
rect 6025 42950 6037 43002
rect 6089 42950 6101 43002
rect 6153 42950 9109 43002
rect 9161 42950 9173 43002
rect 9225 42950 9237 43002
rect 9289 42950 9301 43002
rect 9353 42950 9365 43002
rect 9417 42950 10856 43002
rect 1104 42928 10856 42950
rect 4062 42752 4068 42764
rect 4023 42724 4068 42752
rect 4062 42712 4068 42724
rect 4120 42712 4126 42764
rect 1673 42687 1731 42693
rect 1673 42653 1685 42687
rect 1719 42684 1731 42687
rect 1854 42684 1860 42696
rect 1719 42656 1860 42684
rect 1719 42653 1731 42656
rect 1673 42647 1731 42653
rect 1854 42644 1860 42656
rect 1912 42644 1918 42696
rect 3789 42687 3847 42693
rect 3789 42653 3801 42687
rect 3835 42684 3847 42687
rect 3970 42684 3976 42696
rect 3835 42656 3976 42684
rect 3835 42653 3847 42656
rect 3789 42647 3847 42653
rect 3970 42644 3976 42656
rect 4028 42684 4034 42696
rect 9490 42684 9496 42696
rect 4028 42656 9496 42684
rect 4028 42644 4034 42656
rect 9490 42644 9496 42656
rect 9548 42644 9554 42696
rect 10134 42684 10140 42696
rect 10095 42656 10140 42684
rect 10134 42644 10140 42656
rect 10192 42644 10198 42696
rect 1486 42548 1492 42560
rect 1447 42520 1492 42548
rect 1486 42508 1492 42520
rect 1544 42508 1550 42560
rect 9950 42548 9956 42560
rect 9911 42520 9956 42548
rect 9950 42508 9956 42520
rect 10008 42508 10014 42560
rect 1104 42458 10856 42480
rect 1104 42406 4213 42458
rect 4265 42406 4277 42458
rect 4329 42406 4341 42458
rect 4393 42406 4405 42458
rect 4457 42406 4469 42458
rect 4521 42406 7477 42458
rect 7529 42406 7541 42458
rect 7593 42406 7605 42458
rect 7657 42406 7669 42458
rect 7721 42406 7733 42458
rect 7785 42406 10856 42458
rect 1104 42384 10856 42406
rect 937 42347 995 42353
rect 937 42313 949 42347
rect 983 42344 995 42347
rect 1394 42344 1400 42356
rect 983 42316 1400 42344
rect 983 42313 995 42316
rect 937 42307 995 42313
rect 1394 42304 1400 42316
rect 1452 42304 1458 42356
rect 1394 42168 1400 42220
rect 1452 42208 1458 42220
rect 1673 42211 1731 42217
rect 1673 42208 1685 42211
rect 1452 42180 1685 42208
rect 1452 42168 1458 42180
rect 1673 42177 1685 42180
rect 1719 42177 1731 42211
rect 1673 42171 1731 42177
rect 3973 42211 4031 42217
rect 3973 42177 3985 42211
rect 4019 42208 4031 42211
rect 9858 42208 9864 42220
rect 4019 42180 9864 42208
rect 4019 42177 4031 42180
rect 3973 42171 4031 42177
rect 9858 42168 9864 42180
rect 9916 42168 9922 42220
rect 10134 42208 10140 42220
rect 10095 42180 10140 42208
rect 10134 42168 10140 42180
rect 10192 42168 10198 42220
rect 1486 42004 1492 42016
rect 1447 41976 1492 42004
rect 1486 41964 1492 41976
rect 1544 41964 1550 42016
rect 3970 42004 3976 42016
rect 3931 41976 3976 42004
rect 3970 41964 3976 41976
rect 4028 41964 4034 42016
rect 9858 41964 9864 42016
rect 9916 42004 9922 42016
rect 9953 42007 10011 42013
rect 9953 42004 9965 42007
rect 9916 41976 9965 42004
rect 9916 41964 9922 41976
rect 9953 41973 9965 41976
rect 9999 41973 10011 42007
rect 9953 41967 10011 41973
rect 1104 41914 10856 41936
rect 1104 41862 2582 41914
rect 2634 41862 2646 41914
rect 2698 41862 2710 41914
rect 2762 41862 2774 41914
rect 2826 41862 2838 41914
rect 2890 41862 5845 41914
rect 5897 41862 5909 41914
rect 5961 41862 5973 41914
rect 6025 41862 6037 41914
rect 6089 41862 6101 41914
rect 6153 41862 9109 41914
rect 9161 41862 9173 41914
rect 9225 41862 9237 41914
rect 9289 41862 9301 41914
rect 9353 41862 9365 41914
rect 9417 41862 10856 41914
rect 1104 41840 10856 41862
rect 1302 41760 1308 41812
rect 1360 41800 1366 41812
rect 2133 41803 2191 41809
rect 2133 41800 2145 41803
rect 1360 41772 2145 41800
rect 1360 41760 1366 41772
rect 2133 41769 2145 41772
rect 2179 41769 2191 41803
rect 2133 41763 2191 41769
rect 4062 41732 4068 41744
rect 1688 41704 4068 41732
rect 1688 41605 1716 41704
rect 4062 41692 4068 41704
rect 4120 41692 4126 41744
rect 1673 41599 1731 41605
rect 1673 41565 1685 41599
rect 1719 41565 1731 41599
rect 2130 41596 2136 41608
rect 2091 41568 2136 41596
rect 1673 41559 1731 41565
rect 2130 41556 2136 41568
rect 2188 41556 2194 41608
rect 2317 41599 2375 41605
rect 2317 41565 2329 41599
rect 2363 41596 2375 41599
rect 2774 41596 2780 41608
rect 2363 41568 2780 41596
rect 2363 41565 2375 41568
rect 2317 41559 2375 41565
rect 2774 41556 2780 41568
rect 2832 41596 2838 41608
rect 3510 41596 3516 41608
rect 2832 41568 3516 41596
rect 2832 41556 2838 41568
rect 3510 41556 3516 41568
rect 3568 41556 3574 41608
rect 4065 41599 4123 41605
rect 4065 41565 4077 41599
rect 4111 41596 4123 41599
rect 9766 41596 9772 41608
rect 4111 41568 9772 41596
rect 4111 41565 4123 41568
rect 4065 41559 4123 41565
rect 9766 41556 9772 41568
rect 9824 41556 9830 41608
rect 845 41531 903 41537
rect 845 41497 857 41531
rect 891 41528 903 41531
rect 1302 41528 1308 41540
rect 891 41500 1308 41528
rect 891 41497 903 41500
rect 845 41491 903 41497
rect 1302 41488 1308 41500
rect 1360 41488 1366 41540
rect 2682 41488 2688 41540
rect 2740 41528 2746 41540
rect 3789 41531 3847 41537
rect 3789 41528 3801 41531
rect 2740 41500 3801 41528
rect 2740 41488 2746 41500
rect 3789 41497 3801 41500
rect 3835 41528 3847 41531
rect 4154 41528 4160 41540
rect 3835 41500 4160 41528
rect 3835 41497 3847 41500
rect 3789 41491 3847 41497
rect 4154 41488 4160 41500
rect 4212 41488 4218 41540
rect 1486 41460 1492 41472
rect 1447 41432 1492 41460
rect 1486 41420 1492 41432
rect 1544 41420 1550 41472
rect 1104 41370 10856 41392
rect 1104 41318 4213 41370
rect 4265 41318 4277 41370
rect 4329 41318 4341 41370
rect 4393 41318 4405 41370
rect 4457 41318 4469 41370
rect 4521 41318 7477 41370
rect 7529 41318 7541 41370
rect 7593 41318 7605 41370
rect 7657 41318 7669 41370
rect 7721 41318 7733 41370
rect 7785 41318 10856 41370
rect 1104 41296 10856 41318
rect 1302 41216 1308 41268
rect 1360 41256 1366 41268
rect 1486 41256 1492 41268
rect 1360 41228 1492 41256
rect 1360 41216 1366 41228
rect 1486 41216 1492 41228
rect 1544 41216 1550 41268
rect 1946 41216 1952 41268
rect 2004 41256 2010 41268
rect 2225 41259 2283 41265
rect 2225 41256 2237 41259
rect 2004 41228 2237 41256
rect 2004 41216 2010 41228
rect 2225 41225 2237 41228
rect 2271 41225 2283 41259
rect 2225 41219 2283 41225
rect 3142 41216 3148 41268
rect 3200 41256 3206 41268
rect 3510 41256 3516 41268
rect 3200 41228 3516 41256
rect 3200 41216 3206 41228
rect 3510 41216 3516 41228
rect 3568 41216 3574 41268
rect 2869 41191 2927 41197
rect 2148 41160 2820 41188
rect 2148 41132 2176 41160
rect 1673 41123 1731 41129
rect 1673 41089 1685 41123
rect 1719 41089 1731 41123
rect 2130 41120 2136 41132
rect 2091 41092 2136 41120
rect 1673 41083 1731 41089
rect 1688 40984 1716 41083
rect 2130 41080 2136 41092
rect 2188 41080 2194 41132
rect 2317 41123 2375 41129
rect 2317 41089 2329 41123
rect 2363 41120 2375 41123
rect 2682 41120 2688 41132
rect 2363 41092 2688 41120
rect 2363 41089 2375 41092
rect 2317 41083 2375 41089
rect 2682 41080 2688 41092
rect 2740 41080 2746 41132
rect 2792 41129 2820 41160
rect 2869 41157 2881 41191
rect 2915 41188 2927 41191
rect 3878 41188 3884 41200
rect 2915 41160 3884 41188
rect 2915 41157 2927 41160
rect 2869 41151 2927 41157
rect 3878 41148 3884 41160
rect 3936 41148 3942 41200
rect 6454 41148 6460 41200
rect 6512 41188 6518 41200
rect 6638 41188 6644 41200
rect 6512 41160 6644 41188
rect 6512 41148 6518 41160
rect 6638 41148 6644 41160
rect 6696 41148 6702 41200
rect 2777 41123 2835 41129
rect 2777 41089 2789 41123
rect 2823 41089 2835 41123
rect 2777 41083 2835 41089
rect 2961 41123 3019 41129
rect 2961 41089 2973 41123
rect 3007 41120 3019 41123
rect 3970 41120 3976 41132
rect 3007 41092 3976 41120
rect 3007 41089 3019 41092
rect 2961 41083 3019 41089
rect 3970 41080 3976 41092
rect 4028 41080 4034 41132
rect 4065 41123 4123 41129
rect 4065 41089 4077 41123
rect 4111 41120 4123 41123
rect 9950 41120 9956 41132
rect 4111 41092 9956 41120
rect 4111 41089 4123 41092
rect 4065 41083 4123 41089
rect 9950 41080 9956 41092
rect 10008 41080 10014 41132
rect 10134 41120 10140 41132
rect 10095 41092 10140 41120
rect 10134 41080 10140 41092
rect 10192 41080 10198 41132
rect 3878 40984 3884 40996
rect 1688 40956 3188 40984
rect 1486 40916 1492 40928
rect 1447 40888 1492 40916
rect 1486 40876 1492 40888
rect 1544 40876 1550 40928
rect 3160 40916 3188 40956
rect 3344 40956 3884 40984
rect 3344 40916 3372 40956
rect 3878 40944 3884 40956
rect 3936 40944 3942 40996
rect 3160 40888 3372 40916
rect 4157 40919 4215 40925
rect 4157 40885 4169 40919
rect 4203 40916 4215 40919
rect 4430 40916 4436 40928
rect 4203 40888 4436 40916
rect 4203 40885 4215 40888
rect 4157 40879 4215 40885
rect 4430 40876 4436 40888
rect 4488 40916 4494 40928
rect 6546 40916 6552 40928
rect 4488 40888 6552 40916
rect 4488 40876 4494 40888
rect 6546 40876 6552 40888
rect 6604 40876 6610 40928
rect 9950 40916 9956 40928
rect 9911 40888 9956 40916
rect 9950 40876 9956 40888
rect 10008 40876 10014 40928
rect 1104 40826 10856 40848
rect 1104 40774 2582 40826
rect 2634 40774 2646 40826
rect 2698 40774 2710 40826
rect 2762 40774 2774 40826
rect 2826 40774 2838 40826
rect 2890 40774 5845 40826
rect 5897 40774 5909 40826
rect 5961 40774 5973 40826
rect 6025 40774 6037 40826
rect 6089 40774 6101 40826
rect 6153 40774 9109 40826
rect 9161 40774 9173 40826
rect 9225 40774 9237 40826
rect 9289 40774 9301 40826
rect 9353 40774 9365 40826
rect 9417 40774 10856 40826
rect 1104 40752 10856 40774
rect 1394 40672 1400 40724
rect 1452 40712 1458 40724
rect 2133 40715 2191 40721
rect 2133 40712 2145 40715
rect 1452 40684 2145 40712
rect 1452 40672 1458 40684
rect 2133 40681 2145 40684
rect 2179 40681 2191 40715
rect 2133 40675 2191 40681
rect 2777 40715 2835 40721
rect 2777 40681 2789 40715
rect 2823 40712 2835 40715
rect 3602 40712 3608 40724
rect 2823 40684 3608 40712
rect 2823 40681 2835 40684
rect 2777 40675 2835 40681
rect 3602 40672 3608 40684
rect 3660 40672 3666 40724
rect 3789 40715 3847 40721
rect 3789 40681 3801 40715
rect 3835 40712 3847 40715
rect 4430 40712 4436 40724
rect 3835 40684 4436 40712
rect 3835 40681 3847 40684
rect 3789 40675 3847 40681
rect 4430 40672 4436 40684
rect 4488 40672 4494 40724
rect 2746 40616 4016 40644
rect 2746 40576 2774 40616
rect 2332 40548 2774 40576
rect 1578 40468 1584 40520
rect 1636 40508 1642 40520
rect 1673 40511 1731 40517
rect 1673 40508 1685 40511
rect 1636 40480 1685 40508
rect 1636 40468 1642 40480
rect 1673 40477 1685 40480
rect 1719 40477 1731 40511
rect 2130 40508 2136 40520
rect 2043 40480 2136 40508
rect 1673 40471 1731 40477
rect 2130 40468 2136 40480
rect 2188 40468 2194 40520
rect 2332 40517 2360 40548
rect 2317 40511 2375 40517
rect 2317 40477 2329 40511
rect 2363 40477 2375 40511
rect 2317 40471 2375 40477
rect 2777 40511 2835 40517
rect 2777 40477 2789 40511
rect 2823 40508 2835 40511
rect 2866 40508 2872 40520
rect 2823 40480 2872 40508
rect 2823 40477 2835 40480
rect 2777 40471 2835 40477
rect 2148 40440 2176 40468
rect 2792 40440 2820 40471
rect 2866 40468 2872 40480
rect 2924 40468 2930 40520
rect 2961 40511 3019 40517
rect 2961 40477 2973 40511
rect 3007 40508 3019 40511
rect 3789 40511 3847 40517
rect 3789 40508 3801 40511
rect 3007 40480 3801 40508
rect 3007 40477 3019 40480
rect 2961 40471 3019 40477
rect 3789 40477 3801 40480
rect 3835 40477 3847 40511
rect 3789 40471 3847 40477
rect 2148 40412 2820 40440
rect 1486 40372 1492 40384
rect 1447 40344 1492 40372
rect 1486 40332 1492 40344
rect 1544 40332 1550 40384
rect 3988 40381 4016 40616
rect 4614 40604 4620 40656
rect 4672 40644 4678 40656
rect 5166 40644 5172 40656
rect 4672 40616 5172 40644
rect 4672 40604 4678 40616
rect 5166 40604 5172 40616
rect 5224 40604 5230 40656
rect 5074 40536 5080 40588
rect 5132 40576 5138 40588
rect 5350 40576 5356 40588
rect 5132 40548 5356 40576
rect 5132 40536 5138 40548
rect 5350 40536 5356 40548
rect 5408 40536 5414 40588
rect 4065 40511 4123 40517
rect 4065 40477 4077 40511
rect 4111 40508 4123 40511
rect 9858 40508 9864 40520
rect 4111 40480 9864 40508
rect 4111 40477 4123 40480
rect 4065 40471 4123 40477
rect 9858 40468 9864 40480
rect 9916 40468 9922 40520
rect 10134 40508 10140 40520
rect 10095 40480 10140 40508
rect 10134 40468 10140 40480
rect 10192 40468 10198 40520
rect 3973 40375 4031 40381
rect 3973 40341 3985 40375
rect 4019 40372 4031 40375
rect 6822 40372 6828 40384
rect 4019 40344 6828 40372
rect 4019 40341 4031 40344
rect 3973 40335 4031 40341
rect 6822 40332 6828 40344
rect 6880 40332 6886 40384
rect 9858 40332 9864 40384
rect 9916 40372 9922 40384
rect 9953 40375 10011 40381
rect 9953 40372 9965 40375
rect 9916 40344 9965 40372
rect 9916 40332 9922 40344
rect 9953 40341 9965 40344
rect 9999 40341 10011 40375
rect 9953 40335 10011 40341
rect 1104 40282 10856 40304
rect 1104 40230 4213 40282
rect 4265 40230 4277 40282
rect 4329 40230 4341 40282
rect 4393 40230 4405 40282
rect 4457 40230 4469 40282
rect 4521 40230 7477 40282
rect 7529 40230 7541 40282
rect 7593 40230 7605 40282
rect 7657 40230 7669 40282
rect 7721 40230 7733 40282
rect 7785 40230 10856 40282
rect 1104 40208 10856 40230
rect 3970 40128 3976 40180
rect 4028 40168 4034 40180
rect 5350 40168 5356 40180
rect 4028 40140 5356 40168
rect 4028 40128 4034 40140
rect 5350 40128 5356 40140
rect 5408 40128 5414 40180
rect 9950 40100 9956 40112
rect 4172 40072 9956 40100
rect 1394 40032 1400 40044
rect 1355 40004 1400 40032
rect 1394 39992 1400 40004
rect 1452 39992 1458 40044
rect 2590 40032 2596 40044
rect 2551 40004 2596 40032
rect 2590 39992 2596 40004
rect 2648 39992 2654 40044
rect 2866 40032 2872 40044
rect 2827 40004 2872 40032
rect 2866 39992 2872 40004
rect 2924 39992 2930 40044
rect 4172 40041 4200 40072
rect 9950 40060 9956 40072
rect 10008 40060 10014 40112
rect 4157 40035 4215 40041
rect 4157 40001 4169 40035
rect 4203 40001 4215 40035
rect 10134 40032 10140 40044
rect 10095 40004 10140 40032
rect 4157 39995 4215 40001
rect 10134 39992 10140 40004
rect 10192 39992 10198 40044
rect 1581 39899 1639 39905
rect 1581 39865 1593 39899
rect 1627 39896 1639 39899
rect 5534 39896 5540 39908
rect 1627 39868 5540 39896
rect 1627 39865 1639 39868
rect 1581 39859 1639 39865
rect 5534 39856 5540 39868
rect 5592 39856 5598 39908
rect 3973 39831 4031 39837
rect 3973 39797 3985 39831
rect 4019 39828 4031 39831
rect 5074 39828 5080 39840
rect 4019 39800 5080 39828
rect 4019 39797 4031 39800
rect 3973 39791 4031 39797
rect 5074 39788 5080 39800
rect 5132 39788 5138 39840
rect 9950 39828 9956 39840
rect 9911 39800 9956 39828
rect 9950 39788 9956 39800
rect 10008 39788 10014 39840
rect 1104 39738 10856 39760
rect 1104 39686 2582 39738
rect 2634 39686 2646 39738
rect 2698 39686 2710 39738
rect 2762 39686 2774 39738
rect 2826 39686 2838 39738
rect 2890 39686 5845 39738
rect 5897 39686 5909 39738
rect 5961 39686 5973 39738
rect 6025 39686 6037 39738
rect 6089 39686 6101 39738
rect 6153 39686 9109 39738
rect 9161 39686 9173 39738
rect 9225 39686 9237 39738
rect 9289 39686 9301 39738
rect 9353 39686 9365 39738
rect 9417 39686 10856 39738
rect 1104 39664 10856 39686
rect 2133 39627 2191 39633
rect 2133 39593 2145 39627
rect 2179 39624 2191 39627
rect 2406 39624 2412 39636
rect 2179 39596 2412 39624
rect 2179 39593 2191 39596
rect 2133 39587 2191 39593
rect 2406 39584 2412 39596
rect 2464 39584 2470 39636
rect 1581 39559 1639 39565
rect 1581 39525 1593 39559
rect 1627 39556 1639 39559
rect 5258 39556 5264 39568
rect 1627 39528 5264 39556
rect 1627 39525 1639 39528
rect 1581 39519 1639 39525
rect 5258 39516 5264 39528
rect 5316 39516 5322 39568
rect 937 39491 995 39497
rect 937 39457 949 39491
rect 983 39488 995 39491
rect 2406 39488 2412 39500
rect 983 39460 2412 39488
rect 983 39457 995 39460
rect 937 39451 995 39457
rect 2406 39448 2412 39460
rect 2464 39448 2470 39500
rect 1394 39420 1400 39432
rect 1355 39392 1400 39420
rect 1394 39380 1400 39392
rect 1452 39380 1458 39432
rect 2130 39420 2136 39432
rect 2091 39392 2136 39420
rect 2130 39380 2136 39392
rect 2188 39380 2194 39432
rect 2317 39423 2375 39429
rect 2317 39389 2329 39423
rect 2363 39389 2375 39423
rect 2317 39383 2375 39389
rect 4065 39423 4123 39429
rect 4065 39389 4077 39423
rect 4111 39420 4123 39423
rect 9858 39420 9864 39432
rect 4111 39392 9864 39420
rect 4111 39389 4123 39392
rect 4065 39383 4123 39389
rect 290 39312 296 39364
rect 348 39352 354 39364
rect 2332 39352 2360 39383
rect 9858 39380 9864 39392
rect 9916 39380 9922 39432
rect 3789 39355 3847 39361
rect 3789 39352 3801 39355
rect 348 39324 3801 39352
rect 348 39312 354 39324
rect 3789 39321 3801 39324
rect 3835 39321 3847 39355
rect 3789 39315 3847 39321
rect 1104 39194 10856 39216
rect 1104 39142 4213 39194
rect 4265 39142 4277 39194
rect 4329 39142 4341 39194
rect 4393 39142 4405 39194
rect 4457 39142 4469 39194
rect 4521 39142 7477 39194
rect 7529 39142 7541 39194
rect 7593 39142 7605 39194
rect 7657 39142 7669 39194
rect 7721 39142 7733 39194
rect 7785 39142 10856 39194
rect 1104 39120 10856 39142
rect 1118 39040 1124 39092
rect 1176 39080 1182 39092
rect 1581 39083 1639 39089
rect 1581 39080 1593 39083
rect 1176 39052 1593 39080
rect 1176 39040 1182 39052
rect 1581 39049 1593 39052
rect 1627 39049 1639 39083
rect 1581 39043 1639 39049
rect 1762 39040 1768 39092
rect 1820 39080 1826 39092
rect 2225 39083 2283 39089
rect 2225 39080 2237 39083
rect 1820 39052 2237 39080
rect 1820 39040 1826 39052
rect 2225 39049 2237 39052
rect 2271 39049 2283 39083
rect 2225 39043 2283 39049
rect 2869 39083 2927 39089
rect 2869 39049 2881 39083
rect 2915 39080 2927 39083
rect 3142 39080 3148 39092
rect 2915 39052 3148 39080
rect 2915 39049 2927 39052
rect 2869 39043 2927 39049
rect 3142 39040 3148 39052
rect 3200 39040 3206 39092
rect 2148 38984 2820 39012
rect 2148 38956 2176 38984
rect 1394 38944 1400 38956
rect 1355 38916 1400 38944
rect 1394 38904 1400 38916
rect 1452 38904 1458 38956
rect 2130 38944 2136 38956
rect 2091 38916 2136 38944
rect 2130 38904 2136 38916
rect 2188 38904 2194 38956
rect 2792 38953 2820 38984
rect 2317 38947 2375 38953
rect 2317 38913 2329 38947
rect 2363 38913 2375 38947
rect 2317 38907 2375 38913
rect 2777 38947 2835 38953
rect 2777 38913 2789 38947
rect 2823 38913 2835 38947
rect 2777 38907 2835 38913
rect 2961 38947 3019 38953
rect 2961 38913 2973 38947
rect 3007 38944 3019 38947
rect 5074 38944 5080 38956
rect 3007 38916 5080 38944
rect 3007 38913 3019 38916
rect 2961 38907 3019 38913
rect 1302 38836 1308 38888
rect 1360 38876 1366 38888
rect 1762 38876 1768 38888
rect 1360 38848 1768 38876
rect 1360 38836 1366 38848
rect 1762 38836 1768 38848
rect 1820 38836 1826 38888
rect 2332 38876 2360 38907
rect 5074 38904 5080 38916
rect 5132 38904 5138 38956
rect 10134 38944 10140 38956
rect 10095 38916 10140 38944
rect 10134 38904 10140 38916
rect 10192 38904 10198 38956
rect 3878 38876 3884 38888
rect 2332 38848 3884 38876
rect 3878 38836 3884 38848
rect 3936 38836 3942 38888
rect 9858 38700 9864 38752
rect 9916 38740 9922 38752
rect 9953 38743 10011 38749
rect 9953 38740 9965 38743
rect 9916 38712 9965 38740
rect 9916 38700 9922 38712
rect 9953 38709 9965 38712
rect 9999 38709 10011 38743
rect 9953 38703 10011 38709
rect 1104 38650 10856 38672
rect 1104 38598 2582 38650
rect 2634 38598 2646 38650
rect 2698 38598 2710 38650
rect 2762 38598 2774 38650
rect 2826 38598 2838 38650
rect 2890 38598 5845 38650
rect 5897 38598 5909 38650
rect 5961 38598 5973 38650
rect 6025 38598 6037 38650
rect 6089 38598 6101 38650
rect 6153 38598 9109 38650
rect 9161 38598 9173 38650
rect 9225 38598 9237 38650
rect 9289 38598 9301 38650
rect 9353 38598 9365 38650
rect 9417 38598 10856 38650
rect 1104 38576 10856 38598
rect 2133 38539 2191 38545
rect 2133 38505 2145 38539
rect 2179 38536 2191 38539
rect 2314 38536 2320 38548
rect 2179 38508 2320 38536
rect 2179 38505 2191 38508
rect 2133 38499 2191 38505
rect 2314 38496 2320 38508
rect 2372 38496 2378 38548
rect 2777 38539 2835 38545
rect 2777 38505 2789 38539
rect 2823 38536 2835 38539
rect 3786 38536 3792 38548
rect 2823 38508 3792 38536
rect 2823 38505 2835 38508
rect 2777 38499 2835 38505
rect 3786 38496 3792 38508
rect 3844 38496 3850 38548
rect 1581 38471 1639 38477
rect 1581 38437 1593 38471
rect 1627 38468 1639 38471
rect 7006 38468 7012 38480
rect 1627 38440 7012 38468
rect 1627 38437 1639 38440
rect 1581 38431 1639 38437
rect 7006 38428 7012 38440
rect 7064 38428 7070 38480
rect 1302 38360 1308 38412
rect 1360 38400 1366 38412
rect 1360 38372 2360 38400
rect 1360 38360 1366 38372
rect 1394 38332 1400 38344
rect 1355 38304 1400 38332
rect 1394 38292 1400 38304
rect 1452 38292 1458 38344
rect 2130 38332 2136 38344
rect 2043 38304 2136 38332
rect 2130 38292 2136 38304
rect 2188 38292 2194 38344
rect 2332 38341 2360 38372
rect 2317 38335 2375 38341
rect 2317 38301 2329 38335
rect 2363 38301 2375 38335
rect 2774 38332 2780 38344
rect 2317 38295 2375 38301
rect 2746 38292 2780 38332
rect 2832 38332 2838 38344
rect 2961 38335 3019 38341
rect 2832 38304 2925 38332
rect 2832 38292 2838 38304
rect 2961 38301 2973 38335
rect 3007 38332 3019 38335
rect 4065 38335 4123 38341
rect 3007 38304 3924 38332
rect 3007 38301 3019 38304
rect 2961 38295 3019 38301
rect 2148 38264 2176 38292
rect 2746 38264 2774 38292
rect 2148 38236 2774 38264
rect 750 38156 756 38208
rect 808 38196 814 38208
rect 3602 38196 3608 38208
rect 808 38168 3608 38196
rect 808 38156 814 38168
rect 3602 38156 3608 38168
rect 3660 38156 3666 38208
rect 3896 38205 3924 38304
rect 4065 38301 4077 38335
rect 4111 38332 4123 38335
rect 9950 38332 9956 38344
rect 4111 38304 9956 38332
rect 4111 38301 4123 38304
rect 4065 38295 4123 38301
rect 9950 38292 9956 38304
rect 10008 38292 10014 38344
rect 10134 38332 10140 38344
rect 10095 38304 10140 38332
rect 10134 38292 10140 38304
rect 10192 38292 10198 38344
rect 3881 38199 3939 38205
rect 3881 38165 3893 38199
rect 3927 38196 3939 38199
rect 5626 38196 5632 38208
rect 3927 38168 5632 38196
rect 3927 38165 3939 38168
rect 3881 38159 3939 38165
rect 5626 38156 5632 38168
rect 5684 38156 5690 38208
rect 9950 38196 9956 38208
rect 9911 38168 9956 38196
rect 9950 38156 9956 38168
rect 10008 38156 10014 38208
rect 1104 38106 10856 38128
rect 1104 38054 4213 38106
rect 4265 38054 4277 38106
rect 4329 38054 4341 38106
rect 4393 38054 4405 38106
rect 4457 38054 4469 38106
rect 4521 38054 7477 38106
rect 7529 38054 7541 38106
rect 7593 38054 7605 38106
rect 7657 38054 7669 38106
rect 7721 38054 7733 38106
rect 7785 38054 10856 38106
rect 1104 38032 10856 38054
rect 1581 37995 1639 38001
rect 1581 37961 1593 37995
rect 1627 37992 1639 37995
rect 6178 37992 6184 38004
rect 1627 37964 6184 37992
rect 1627 37961 1639 37964
rect 1581 37955 1639 37961
rect 6178 37952 6184 37964
rect 6236 37952 6242 38004
rect 1394 37856 1400 37868
rect 1355 37828 1400 37856
rect 1394 37816 1400 37828
rect 1452 37816 1458 37868
rect 2685 37859 2743 37865
rect 2685 37825 2697 37859
rect 2731 37856 2743 37859
rect 2774 37856 2780 37868
rect 2731 37828 2780 37856
rect 2731 37825 2743 37828
rect 2685 37819 2743 37825
rect 2774 37816 2780 37828
rect 2832 37816 2838 37868
rect 3973 37859 4031 37865
rect 3973 37825 3985 37859
rect 4019 37856 4031 37859
rect 9858 37856 9864 37868
rect 4019 37828 9864 37856
rect 4019 37825 4031 37828
rect 3973 37819 4031 37825
rect 9858 37816 9864 37828
rect 9916 37816 9922 37868
rect 2314 37748 2320 37800
rect 2372 37788 2378 37800
rect 2409 37791 2467 37797
rect 2409 37788 2421 37791
rect 2372 37760 2421 37788
rect 2372 37748 2378 37760
rect 2409 37757 2421 37760
rect 2455 37788 2467 37791
rect 3050 37788 3056 37800
rect 2455 37760 3056 37788
rect 2455 37757 2467 37760
rect 2409 37751 2467 37757
rect 3050 37748 3056 37760
rect 3108 37748 3114 37800
rect 3878 37612 3884 37664
rect 3936 37652 3942 37664
rect 3973 37655 4031 37661
rect 3973 37652 3985 37655
rect 3936 37624 3985 37652
rect 3936 37612 3942 37624
rect 3973 37621 3985 37624
rect 4019 37652 4031 37655
rect 6178 37652 6184 37664
rect 4019 37624 6184 37652
rect 4019 37621 4031 37624
rect 3973 37615 4031 37621
rect 6178 37612 6184 37624
rect 6236 37612 6242 37664
rect 1104 37562 10856 37584
rect 1104 37510 2582 37562
rect 2634 37510 2646 37562
rect 2698 37510 2710 37562
rect 2762 37510 2774 37562
rect 2826 37510 2838 37562
rect 2890 37510 5845 37562
rect 5897 37510 5909 37562
rect 5961 37510 5973 37562
rect 6025 37510 6037 37562
rect 6089 37510 6101 37562
rect 6153 37510 9109 37562
rect 9161 37510 9173 37562
rect 9225 37510 9237 37562
rect 9289 37510 9301 37562
rect 9353 37510 9365 37562
rect 9417 37510 10856 37562
rect 1104 37488 10856 37510
rect 382 37340 388 37392
rect 440 37380 446 37392
rect 1302 37380 1308 37392
rect 440 37352 1308 37380
rect 440 37340 446 37352
rect 1302 37340 1308 37352
rect 1360 37380 1366 37392
rect 3881 37383 3939 37389
rect 3881 37380 3893 37383
rect 1360 37352 3893 37380
rect 1360 37340 1366 37352
rect 3881 37349 3893 37352
rect 3927 37349 3939 37383
rect 3881 37343 3939 37349
rect 2314 37272 2320 37324
rect 2372 37312 2378 37324
rect 2409 37315 2467 37321
rect 2409 37312 2421 37315
rect 2372 37284 2421 37312
rect 2372 37272 2378 37284
rect 2409 37281 2421 37284
rect 2455 37281 2467 37315
rect 2409 37275 2467 37281
rect 1394 37244 1400 37256
rect 1355 37216 1400 37244
rect 1394 37204 1400 37216
rect 1452 37204 1458 37256
rect 2682 37244 2688 37256
rect 2643 37216 2688 37244
rect 2682 37204 2688 37216
rect 2740 37204 2746 37256
rect 4065 37247 4123 37253
rect 4065 37213 4077 37247
rect 4111 37244 4123 37247
rect 9950 37244 9956 37256
rect 4111 37216 9956 37244
rect 4111 37213 4123 37216
rect 4065 37207 4123 37213
rect 9950 37204 9956 37216
rect 10008 37204 10014 37256
rect 10134 37244 10140 37256
rect 10095 37216 10140 37244
rect 10134 37204 10140 37216
rect 10192 37204 10198 37256
rect 3050 37136 3056 37188
rect 3108 37176 3114 37188
rect 4982 37176 4988 37188
rect 3108 37148 4988 37176
rect 3108 37136 3114 37148
rect 4982 37136 4988 37148
rect 5040 37136 5046 37188
rect 1581 37111 1639 37117
rect 1581 37077 1593 37111
rect 1627 37108 1639 37111
rect 6454 37108 6460 37120
rect 1627 37080 6460 37108
rect 1627 37077 1639 37080
rect 1581 37071 1639 37077
rect 6454 37068 6460 37080
rect 6512 37068 6518 37120
rect 9950 37108 9956 37120
rect 9911 37080 9956 37108
rect 9950 37068 9956 37080
rect 10008 37068 10014 37120
rect 1104 37018 10856 37040
rect 1104 36966 4213 37018
rect 4265 36966 4277 37018
rect 4329 36966 4341 37018
rect 4393 36966 4405 37018
rect 4457 36966 4469 37018
rect 4521 36966 7477 37018
rect 7529 36966 7541 37018
rect 7593 36966 7605 37018
rect 7657 36966 7669 37018
rect 7721 36966 7733 37018
rect 7785 36966 10856 37018
rect 1104 36944 10856 36966
rect 1946 36864 1952 36916
rect 2004 36904 2010 36916
rect 2225 36907 2283 36913
rect 2225 36904 2237 36907
rect 2004 36876 2237 36904
rect 2004 36864 2010 36876
rect 2225 36873 2237 36876
rect 2271 36873 2283 36907
rect 2225 36867 2283 36873
rect 2869 36907 2927 36913
rect 2869 36873 2881 36907
rect 2915 36904 2927 36907
rect 3694 36904 3700 36916
rect 2915 36876 3700 36904
rect 2915 36873 2927 36876
rect 2869 36867 2927 36873
rect 3694 36864 3700 36876
rect 3752 36864 3758 36916
rect 2682 36836 2688 36848
rect 2148 36808 2688 36836
rect 2148 36780 2176 36808
rect 2682 36796 2688 36808
rect 2740 36836 2746 36848
rect 3786 36836 3792 36848
rect 2740 36808 2820 36836
rect 2740 36796 2746 36808
rect 1394 36768 1400 36780
rect 1355 36740 1400 36768
rect 1394 36728 1400 36740
rect 1452 36728 1458 36780
rect 2130 36768 2136 36780
rect 2043 36740 2136 36768
rect 2130 36728 2136 36740
rect 2188 36728 2194 36780
rect 2792 36777 2820 36808
rect 2884 36808 3792 36836
rect 2317 36771 2375 36777
rect 2317 36737 2329 36771
rect 2363 36737 2375 36771
rect 2317 36731 2375 36737
rect 2777 36771 2835 36777
rect 2777 36737 2789 36771
rect 2823 36737 2835 36771
rect 2777 36731 2835 36737
rect 1118 36660 1124 36712
rect 1176 36700 1182 36712
rect 2332 36700 2360 36731
rect 2884 36700 2912 36808
rect 3786 36796 3792 36808
rect 3844 36796 3850 36848
rect 2961 36771 3019 36777
rect 2961 36737 2973 36771
rect 3007 36768 3019 36771
rect 4065 36771 4123 36777
rect 4065 36768 4077 36771
rect 3007 36740 4077 36768
rect 3007 36737 3019 36740
rect 2961 36731 3019 36737
rect 4065 36737 4077 36740
rect 4111 36737 4123 36771
rect 4065 36731 4123 36737
rect 4341 36771 4399 36777
rect 4341 36737 4353 36771
rect 4387 36768 4399 36771
rect 9950 36768 9956 36780
rect 4387 36740 9956 36768
rect 4387 36737 4399 36740
rect 4341 36731 4399 36737
rect 1176 36672 2268 36700
rect 2332 36672 2912 36700
rect 1176 36660 1182 36672
rect 2240 36632 2268 36672
rect 2976 36632 3004 36731
rect 9950 36728 9956 36740
rect 10008 36728 10014 36780
rect 10134 36768 10140 36780
rect 10095 36740 10140 36768
rect 10134 36728 10140 36740
rect 10192 36728 10198 36780
rect 4798 36632 4804 36644
rect 2240 36604 3004 36632
rect 3252 36604 4804 36632
rect 14 36524 20 36576
rect 72 36564 78 36576
rect 750 36564 756 36576
rect 72 36536 756 36564
rect 72 36524 78 36536
rect 750 36524 756 36536
rect 808 36524 814 36576
rect 1581 36567 1639 36573
rect 1581 36533 1593 36567
rect 1627 36564 1639 36567
rect 3252 36564 3280 36604
rect 4798 36592 4804 36604
rect 4856 36592 4862 36644
rect 1627 36536 3280 36564
rect 1627 36533 1639 36536
rect 1581 36527 1639 36533
rect 3326 36524 3332 36576
rect 3384 36564 3390 36576
rect 3510 36564 3516 36576
rect 3384 36536 3516 36564
rect 3384 36524 3390 36536
rect 3510 36524 3516 36536
rect 3568 36524 3574 36576
rect 3878 36524 3884 36576
rect 3936 36564 3942 36576
rect 4062 36564 4068 36576
rect 3936 36536 4068 36564
rect 3936 36524 3942 36536
rect 4062 36524 4068 36536
rect 4120 36524 4126 36576
rect 4338 36524 4344 36576
rect 4396 36564 4402 36576
rect 9953 36567 10011 36573
rect 9953 36564 9965 36567
rect 4396 36536 9965 36564
rect 4396 36524 4402 36536
rect 9953 36533 9965 36536
rect 9999 36533 10011 36567
rect 9953 36527 10011 36533
rect 1104 36474 10856 36496
rect 1104 36422 2582 36474
rect 2634 36422 2646 36474
rect 2698 36422 2710 36474
rect 2762 36422 2774 36474
rect 2826 36422 2838 36474
rect 2890 36422 5845 36474
rect 5897 36422 5909 36474
rect 5961 36422 5973 36474
rect 6025 36422 6037 36474
rect 6089 36422 6101 36474
rect 6153 36422 9109 36474
rect 9161 36422 9173 36474
rect 9225 36422 9237 36474
rect 9289 36422 9301 36474
rect 9353 36422 9365 36474
rect 9417 36422 10856 36474
rect 1104 36400 10856 36422
rect 474 36320 480 36372
rect 532 36360 538 36372
rect 1581 36363 1639 36369
rect 1581 36360 1593 36363
rect 532 36332 1593 36360
rect 532 36320 538 36332
rect 1581 36329 1593 36332
rect 1627 36329 1639 36363
rect 1581 36323 1639 36329
rect 2777 36363 2835 36369
rect 2777 36329 2789 36363
rect 2823 36360 2835 36363
rect 3602 36360 3608 36372
rect 2823 36332 3608 36360
rect 2823 36329 2835 36332
rect 2777 36323 2835 36329
rect 3602 36320 3608 36332
rect 3660 36320 3666 36372
rect 1486 36252 1492 36304
rect 1544 36292 1550 36304
rect 2133 36295 2191 36301
rect 2133 36292 2145 36295
rect 1544 36264 2145 36292
rect 1544 36252 1550 36264
rect 2133 36261 2145 36264
rect 2179 36261 2191 36295
rect 2133 36255 2191 36261
rect 4982 36224 4988 36236
rect 2332 36196 4988 36224
rect 1394 36156 1400 36168
rect 1355 36128 1400 36156
rect 1394 36116 1400 36128
rect 1452 36116 1458 36168
rect 2130 36156 2136 36168
rect 2091 36128 2136 36156
rect 2130 36116 2136 36128
rect 2188 36116 2194 36168
rect 2332 36165 2360 36196
rect 4982 36184 4988 36196
rect 5040 36184 5046 36236
rect 2317 36159 2375 36165
rect 2317 36125 2329 36159
rect 2363 36125 2375 36159
rect 2317 36119 2375 36125
rect 2777 36159 2835 36165
rect 2777 36125 2789 36159
rect 2823 36125 2835 36159
rect 2777 36119 2835 36125
rect 2961 36159 3019 36165
rect 2961 36125 2973 36159
rect 3007 36125 3019 36159
rect 2961 36119 3019 36125
rect 2148 36088 2176 36116
rect 2792 36088 2820 36119
rect 2148 36060 2820 36088
rect 2976 36088 3004 36119
rect 3786 36116 3792 36168
rect 3844 36156 3850 36168
rect 4065 36159 4123 36165
rect 4065 36156 4077 36159
rect 3844 36128 4077 36156
rect 3844 36116 3850 36128
rect 4065 36125 4077 36128
rect 4111 36125 4123 36159
rect 4338 36156 4344 36168
rect 4299 36128 4344 36156
rect 4065 36119 4123 36125
rect 4338 36116 4344 36128
rect 4396 36116 4402 36168
rect 10134 36156 10140 36168
rect 10095 36128 10140 36156
rect 10134 36116 10140 36128
rect 10192 36116 10198 36168
rect 4798 36088 4804 36100
rect 2976 36060 4804 36088
rect 4798 36048 4804 36060
rect 4856 36048 4862 36100
rect 1578 35980 1584 36032
rect 1636 36020 1642 36032
rect 5166 36020 5172 36032
rect 1636 35992 5172 36020
rect 1636 35980 1642 35992
rect 5166 35980 5172 35992
rect 5224 35980 5230 36032
rect 9950 36020 9956 36032
rect 9911 35992 9956 36020
rect 9950 35980 9956 35992
rect 10008 35980 10014 36032
rect 1104 35930 10856 35952
rect 1104 35878 4213 35930
rect 4265 35878 4277 35930
rect 4329 35878 4341 35930
rect 4393 35878 4405 35930
rect 4457 35878 4469 35930
rect 4521 35878 7477 35930
rect 7529 35878 7541 35930
rect 7593 35878 7605 35930
rect 7657 35878 7669 35930
rect 7721 35878 7733 35930
rect 7785 35878 10856 35930
rect 1104 35856 10856 35878
rect 1670 35776 1676 35828
rect 1728 35816 1734 35828
rect 2225 35819 2283 35825
rect 2225 35816 2237 35819
rect 1728 35788 2237 35816
rect 1728 35776 1734 35788
rect 2225 35785 2237 35788
rect 2271 35785 2283 35819
rect 5258 35816 5264 35828
rect 2225 35779 2283 35785
rect 4264 35788 5264 35816
rect 4264 35760 4292 35788
rect 5258 35776 5264 35788
rect 5316 35776 5322 35828
rect 4246 35708 4252 35760
rect 4304 35708 4310 35760
rect 1394 35680 1400 35692
rect 1355 35652 1400 35680
rect 1394 35640 1400 35652
rect 1452 35640 1458 35692
rect 2130 35680 2136 35692
rect 2091 35652 2136 35680
rect 2130 35640 2136 35652
rect 2188 35640 2194 35692
rect 2317 35683 2375 35689
rect 2317 35649 2329 35683
rect 2363 35649 2375 35683
rect 2317 35643 2375 35649
rect 4341 35683 4399 35689
rect 4341 35649 4353 35683
rect 4387 35680 4399 35683
rect 9950 35680 9956 35692
rect 4387 35652 9956 35680
rect 4387 35649 4399 35652
rect 4341 35643 4399 35649
rect 474 35572 480 35624
rect 532 35612 538 35624
rect 2332 35612 2360 35643
rect 9950 35640 9956 35652
rect 10008 35640 10014 35692
rect 4065 35615 4123 35621
rect 4065 35612 4077 35615
rect 532 35584 4077 35612
rect 532 35572 538 35584
rect 4065 35581 4077 35584
rect 4111 35581 4123 35615
rect 4065 35575 4123 35581
rect 4614 35572 4620 35624
rect 4672 35612 4678 35624
rect 5442 35612 5448 35624
rect 4672 35584 5448 35612
rect 4672 35572 4678 35584
rect 5442 35572 5448 35584
rect 5500 35572 5506 35624
rect 1581 35547 1639 35553
rect 1581 35513 1593 35547
rect 1627 35544 1639 35547
rect 5534 35544 5540 35556
rect 1627 35516 5540 35544
rect 1627 35513 1639 35516
rect 1581 35507 1639 35513
rect 5534 35504 5540 35516
rect 5592 35504 5598 35556
rect 5166 35436 5172 35488
rect 5224 35476 5230 35488
rect 5350 35476 5356 35488
rect 5224 35448 5356 35476
rect 5224 35436 5230 35448
rect 5350 35436 5356 35448
rect 5408 35436 5414 35488
rect 1104 35386 10856 35408
rect 1104 35334 2582 35386
rect 2634 35334 2646 35386
rect 2698 35334 2710 35386
rect 2762 35334 2774 35386
rect 2826 35334 2838 35386
rect 2890 35334 5845 35386
rect 5897 35334 5909 35386
rect 5961 35334 5973 35386
rect 6025 35334 6037 35386
rect 6089 35334 6101 35386
rect 6153 35334 9109 35386
rect 9161 35334 9173 35386
rect 9225 35334 9237 35386
rect 9289 35334 9301 35386
rect 9353 35334 9365 35386
rect 9417 35334 10856 35386
rect 1104 35312 10856 35334
rect 1210 35232 1216 35284
rect 1268 35272 1274 35284
rect 1581 35275 1639 35281
rect 1581 35272 1593 35275
rect 1268 35244 1593 35272
rect 1268 35232 1274 35244
rect 1581 35241 1593 35244
rect 1627 35241 1639 35275
rect 1581 35235 1639 35241
rect 198 35164 204 35216
rect 256 35204 262 35216
rect 3970 35204 3976 35216
rect 256 35176 3976 35204
rect 256 35164 262 35176
rect 3970 35164 3976 35176
rect 4028 35164 4034 35216
rect 1394 35068 1400 35080
rect 1355 35040 1400 35068
rect 1394 35028 1400 35040
rect 1452 35028 1458 35080
rect 4341 35071 4399 35077
rect 4341 35037 4353 35071
rect 4387 35068 4399 35071
rect 10134 35068 10140 35080
rect 4387 35040 9996 35068
rect 10095 35040 10140 35068
rect 4387 35037 4399 35040
rect 4341 35031 4399 35037
rect 1762 34960 1768 35012
rect 1820 35000 1826 35012
rect 4246 35000 4252 35012
rect 1820 34972 4252 35000
rect 1820 34960 1826 34972
rect 4246 34960 4252 34972
rect 4304 34960 4310 35012
rect 4157 34935 4215 34941
rect 4157 34901 4169 34935
rect 4203 34932 4215 34935
rect 4798 34932 4804 34944
rect 4203 34904 4804 34932
rect 4203 34901 4215 34904
rect 4157 34895 4215 34901
rect 4798 34892 4804 34904
rect 4856 34892 4862 34944
rect 9968 34941 9996 35040
rect 10134 35028 10140 35040
rect 10192 35028 10198 35080
rect 9953 34935 10011 34941
rect 9953 34901 9965 34935
rect 9999 34901 10011 34935
rect 9953 34895 10011 34901
rect 1104 34842 10856 34864
rect 1104 34790 4213 34842
rect 4265 34790 4277 34842
rect 4329 34790 4341 34842
rect 4393 34790 4405 34842
rect 4457 34790 4469 34842
rect 4521 34790 7477 34842
rect 7529 34790 7541 34842
rect 7593 34790 7605 34842
rect 7657 34790 7669 34842
rect 7721 34790 7733 34842
rect 7785 34790 10856 34842
rect 1104 34768 10856 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 4157 34731 4215 34737
rect 1627 34700 2774 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 2746 34660 2774 34700
rect 4157 34697 4169 34731
rect 4203 34728 4215 34731
rect 4982 34728 4988 34740
rect 4203 34700 4988 34728
rect 4203 34697 4215 34700
rect 4157 34691 4215 34697
rect 4982 34688 4988 34700
rect 5040 34728 5046 34740
rect 5350 34728 5356 34740
rect 5040 34700 5356 34728
rect 5040 34688 5046 34700
rect 5350 34688 5356 34700
rect 5408 34688 5414 34740
rect 9953 34731 10011 34737
rect 9953 34697 9965 34731
rect 9999 34697 10011 34731
rect 9953 34691 10011 34697
rect 6638 34660 6644 34672
rect 2746 34632 6644 34660
rect 6638 34620 6644 34632
rect 6696 34620 6702 34672
rect 1394 34592 1400 34604
rect 1355 34564 1400 34592
rect 1394 34552 1400 34564
rect 1452 34552 1458 34604
rect 4341 34595 4399 34601
rect 4341 34561 4353 34595
rect 4387 34592 4399 34595
rect 9968 34592 9996 34691
rect 4387 34564 9996 34592
rect 10137 34595 10195 34601
rect 4387 34561 4399 34564
rect 4341 34555 4399 34561
rect 10137 34561 10149 34595
rect 10183 34561 10195 34595
rect 10137 34555 10195 34561
rect 3786 34484 3792 34536
rect 3844 34524 3850 34536
rect 4982 34524 4988 34536
rect 3844 34496 4988 34524
rect 3844 34484 3850 34496
rect 4982 34484 4988 34496
rect 5040 34484 5046 34536
rect 10152 34468 10180 34555
rect 10134 34416 10140 34468
rect 10192 34416 10198 34468
rect 1104 34298 10856 34320
rect 1104 34246 2582 34298
rect 2634 34246 2646 34298
rect 2698 34246 2710 34298
rect 2762 34246 2774 34298
rect 2826 34246 2838 34298
rect 2890 34246 5845 34298
rect 5897 34246 5909 34298
rect 5961 34246 5973 34298
rect 6025 34246 6037 34298
rect 6089 34246 6101 34298
rect 6153 34246 9109 34298
rect 9161 34246 9173 34298
rect 9225 34246 9237 34298
rect 9289 34246 9301 34298
rect 9353 34246 9365 34298
rect 9417 34246 10856 34298
rect 1104 34224 10856 34246
rect 1581 34187 1639 34193
rect 1581 34153 1593 34187
rect 1627 34184 1639 34187
rect 5718 34184 5724 34196
rect 1627 34156 5724 34184
rect 1627 34153 1639 34156
rect 1581 34147 1639 34153
rect 5718 34144 5724 34156
rect 5776 34144 5782 34196
rect 1394 33980 1400 33992
rect 1355 33952 1400 33980
rect 1394 33940 1400 33952
rect 1452 33940 1458 33992
rect 10134 33980 10140 33992
rect 10095 33952 10140 33980
rect 10134 33940 10140 33952
rect 10192 33940 10198 33992
rect 9858 33804 9864 33856
rect 9916 33844 9922 33856
rect 9953 33847 10011 33853
rect 9953 33844 9965 33847
rect 9916 33816 9965 33844
rect 9916 33804 9922 33816
rect 9953 33813 9965 33816
rect 9999 33813 10011 33847
rect 9953 33807 10011 33813
rect 1104 33754 10856 33776
rect 1104 33702 4213 33754
rect 4265 33702 4277 33754
rect 4329 33702 4341 33754
rect 4393 33702 4405 33754
rect 4457 33702 4469 33754
rect 4521 33702 7477 33754
rect 7529 33702 7541 33754
rect 7593 33702 7605 33754
rect 7657 33702 7669 33754
rect 7721 33702 7733 33754
rect 7785 33702 10856 33754
rect 1104 33680 10856 33702
rect 1578 33640 1584 33652
rect 1539 33612 1584 33640
rect 1578 33600 1584 33612
rect 1636 33600 1642 33652
rect 1394 33504 1400 33516
rect 1355 33476 1400 33504
rect 1394 33464 1400 33476
rect 1452 33464 1458 33516
rect 1104 33210 10856 33232
rect 1104 33158 2582 33210
rect 2634 33158 2646 33210
rect 2698 33158 2710 33210
rect 2762 33158 2774 33210
rect 2826 33158 2838 33210
rect 2890 33158 5845 33210
rect 5897 33158 5909 33210
rect 5961 33158 5973 33210
rect 6025 33158 6037 33210
rect 6089 33158 6101 33210
rect 6153 33158 9109 33210
rect 9161 33158 9173 33210
rect 9225 33158 9237 33210
rect 9289 33158 9301 33210
rect 9353 33158 9365 33210
rect 9417 33158 10856 33210
rect 1104 33136 10856 33158
rect 934 33056 940 33108
rect 992 33096 998 33108
rect 1581 33099 1639 33105
rect 1581 33096 1593 33099
rect 992 33068 1593 33096
rect 992 33056 998 33068
rect 1581 33065 1593 33068
rect 1627 33065 1639 33099
rect 1581 33059 1639 33065
rect 1394 32892 1400 32904
rect 1355 32864 1400 32892
rect 1394 32852 1400 32864
rect 1452 32852 1458 32904
rect 10134 32892 10140 32904
rect 10095 32864 10140 32892
rect 10134 32852 10140 32864
rect 10192 32852 10198 32904
rect 9950 32756 9956 32768
rect 9911 32728 9956 32756
rect 9950 32716 9956 32728
rect 10008 32716 10014 32768
rect 1104 32666 10856 32688
rect 1104 32614 4213 32666
rect 4265 32614 4277 32666
rect 4329 32614 4341 32666
rect 4393 32614 4405 32666
rect 4457 32614 4469 32666
rect 4521 32614 7477 32666
rect 7529 32614 7541 32666
rect 7593 32614 7605 32666
rect 7657 32614 7669 32666
rect 7721 32614 7733 32666
rect 7785 32614 10856 32666
rect 1104 32592 10856 32614
rect 1026 32512 1032 32564
rect 1084 32552 1090 32564
rect 1581 32555 1639 32561
rect 1581 32552 1593 32555
rect 1084 32524 1593 32552
rect 1084 32512 1090 32524
rect 1581 32521 1593 32524
rect 1627 32521 1639 32555
rect 2222 32552 2228 32564
rect 2183 32524 2228 32552
rect 1581 32515 1639 32521
rect 2222 32512 2228 32524
rect 2280 32512 2286 32564
rect 1302 32376 1308 32428
rect 1360 32416 1366 32428
rect 1397 32419 1455 32425
rect 1397 32416 1409 32419
rect 1360 32388 1409 32416
rect 1360 32376 1366 32388
rect 1397 32385 1409 32388
rect 1443 32385 1455 32419
rect 2130 32416 2136 32428
rect 2091 32388 2136 32416
rect 1397 32379 1455 32385
rect 2130 32376 2136 32388
rect 2188 32376 2194 32428
rect 2317 32419 2375 32425
rect 2317 32385 2329 32419
rect 2363 32416 2375 32419
rect 3142 32416 3148 32428
rect 2363 32388 3148 32416
rect 2363 32385 2375 32388
rect 2317 32379 2375 32385
rect 3142 32376 3148 32388
rect 3200 32376 3206 32428
rect 10134 32416 10140 32428
rect 10095 32388 10140 32416
rect 10134 32376 10140 32388
rect 10192 32376 10198 32428
rect 1670 32240 1676 32292
rect 1728 32280 1734 32292
rect 6454 32280 6460 32292
rect 1728 32252 6460 32280
rect 1728 32240 1734 32252
rect 6454 32240 6460 32252
rect 6512 32240 6518 32292
rect 9766 32172 9772 32224
rect 9824 32212 9830 32224
rect 9953 32215 10011 32221
rect 9953 32212 9965 32215
rect 9824 32184 9965 32212
rect 9824 32172 9830 32184
rect 9953 32181 9965 32184
rect 9999 32181 10011 32215
rect 9953 32175 10011 32181
rect 1104 32122 10856 32144
rect 1104 32070 2582 32122
rect 2634 32070 2646 32122
rect 2698 32070 2710 32122
rect 2762 32070 2774 32122
rect 2826 32070 2838 32122
rect 2890 32070 5845 32122
rect 5897 32070 5909 32122
rect 5961 32070 5973 32122
rect 6025 32070 6037 32122
rect 6089 32070 6101 32122
rect 6153 32070 9109 32122
rect 9161 32070 9173 32122
rect 9225 32070 9237 32122
rect 9289 32070 9301 32122
rect 9353 32070 9365 32122
rect 9417 32070 10856 32122
rect 1104 32048 10856 32070
rect 2133 32011 2191 32017
rect 2133 31977 2145 32011
rect 2179 32008 2191 32011
rect 2406 32008 2412 32020
rect 2179 31980 2412 32008
rect 2179 31977 2191 31980
rect 2133 31971 2191 31977
rect 2406 31968 2412 31980
rect 2464 31968 2470 32020
rect 10965 32011 11023 32017
rect 10965 32008 10977 32011
rect 2746 31980 10977 32008
rect 1581 31943 1639 31949
rect 1581 31909 1593 31943
rect 1627 31940 1639 31943
rect 2746 31940 2774 31980
rect 10965 31977 10977 31980
rect 11011 31977 11023 32011
rect 10965 31971 11023 31977
rect 1627 31912 2774 31940
rect 1627 31909 1639 31912
rect 1581 31903 1639 31909
rect 3142 31900 3148 31952
rect 3200 31940 3206 31952
rect 3237 31943 3295 31949
rect 3237 31940 3249 31943
rect 3200 31912 3249 31940
rect 3200 31900 3206 31912
rect 3237 31909 3249 31912
rect 3283 31940 3295 31943
rect 5534 31940 5540 31952
rect 3283 31912 5540 31940
rect 3283 31909 3295 31912
rect 3237 31903 3295 31909
rect 5534 31900 5540 31912
rect 5592 31900 5598 31952
rect 1394 31804 1400 31816
rect 1355 31776 1400 31804
rect 1394 31764 1400 31776
rect 1452 31764 1458 31816
rect 2130 31804 2136 31816
rect 2091 31776 2136 31804
rect 2130 31764 2136 31776
rect 2188 31764 2194 31816
rect 2311 31807 2369 31813
rect 2311 31773 2323 31807
rect 2357 31773 2369 31807
rect 2311 31767 2369 31773
rect 3237 31807 3295 31813
rect 3237 31773 3249 31807
rect 3283 31804 3295 31807
rect 9858 31804 9864 31816
rect 3283 31776 9864 31804
rect 3283 31773 3295 31776
rect 3237 31767 3295 31773
rect 198 31696 204 31748
rect 256 31736 262 31748
rect 2332 31736 2360 31767
rect 9858 31764 9864 31776
rect 9916 31764 9922 31816
rect 3142 31736 3148 31748
rect 256 31708 3148 31736
rect 256 31696 262 31708
rect 3142 31696 3148 31708
rect 3200 31696 3206 31748
rect 1104 31578 10856 31600
rect 1104 31526 4213 31578
rect 4265 31526 4277 31578
rect 4329 31526 4341 31578
rect 4393 31526 4405 31578
rect 4457 31526 4469 31578
rect 4521 31526 7477 31578
rect 7529 31526 7541 31578
rect 7593 31526 7605 31578
rect 7657 31526 7669 31578
rect 7721 31526 7733 31578
rect 7785 31526 10856 31578
rect 1104 31504 10856 31526
rect 1581 31467 1639 31473
rect 1581 31433 1593 31467
rect 1627 31464 1639 31467
rect 1670 31464 1676 31476
rect 1627 31436 1676 31464
rect 1627 31433 1639 31436
rect 1581 31427 1639 31433
rect 1670 31424 1676 31436
rect 1728 31424 1734 31476
rect 2038 31424 2044 31476
rect 2096 31464 2102 31476
rect 2225 31467 2283 31473
rect 2225 31464 2237 31467
rect 2096 31436 2237 31464
rect 2096 31424 2102 31436
rect 2225 31433 2237 31436
rect 2271 31433 2283 31467
rect 3142 31464 3148 31476
rect 3103 31436 3148 31464
rect 2225 31427 2283 31433
rect 3142 31424 3148 31436
rect 3200 31424 3206 31476
rect 1302 31288 1308 31340
rect 1360 31328 1366 31340
rect 1397 31331 1455 31337
rect 1397 31328 1409 31331
rect 1360 31300 1409 31328
rect 1360 31288 1366 31300
rect 1397 31297 1409 31300
rect 1443 31297 1455 31331
rect 2130 31328 2136 31340
rect 2091 31300 2136 31328
rect 1397 31291 1455 31297
rect 2130 31288 2136 31300
rect 2188 31288 2194 31340
rect 2317 31331 2375 31337
rect 2317 31297 2329 31331
rect 2363 31328 2375 31331
rect 3142 31328 3148 31340
rect 2363 31300 3148 31328
rect 2363 31297 2375 31300
rect 2317 31291 2375 31297
rect 3142 31288 3148 31300
rect 3200 31288 3206 31340
rect 3329 31331 3387 31337
rect 3329 31297 3341 31331
rect 3375 31328 3387 31331
rect 9950 31328 9956 31340
rect 3375 31300 9956 31328
rect 3375 31297 3387 31300
rect 3329 31291 3387 31297
rect 9950 31288 9956 31300
rect 10008 31288 10014 31340
rect 10134 31328 10140 31340
rect 10095 31300 10140 31328
rect 10134 31288 10140 31300
rect 10192 31288 10198 31340
rect 1670 31152 1676 31204
rect 1728 31192 1734 31204
rect 8386 31192 8392 31204
rect 1728 31164 8392 31192
rect 1728 31152 1734 31164
rect 8386 31152 8392 31164
rect 8444 31152 8450 31204
rect 3326 31084 3332 31136
rect 3384 31124 3390 31136
rect 4706 31124 4712 31136
rect 3384 31096 4712 31124
rect 3384 31084 3390 31096
rect 4706 31084 4712 31096
rect 4764 31084 4770 31136
rect 9858 31084 9864 31136
rect 9916 31124 9922 31136
rect 9953 31127 10011 31133
rect 9953 31124 9965 31127
rect 9916 31096 9965 31124
rect 9916 31084 9922 31096
rect 9953 31093 9965 31096
rect 9999 31093 10011 31127
rect 9953 31087 10011 31093
rect 1104 31034 10856 31056
rect 1104 30982 2582 31034
rect 2634 30982 2646 31034
rect 2698 30982 2710 31034
rect 2762 30982 2774 31034
rect 2826 30982 2838 31034
rect 2890 30982 5845 31034
rect 5897 30982 5909 31034
rect 5961 30982 5973 31034
rect 6025 30982 6037 31034
rect 6089 30982 6101 31034
rect 6153 30982 9109 31034
rect 9161 30982 9173 31034
rect 9225 30982 9237 31034
rect 9289 30982 9301 31034
rect 9353 30982 9365 31034
rect 9417 30982 10856 31034
rect 1104 30960 10856 30982
rect 1581 30923 1639 30929
rect 1581 30889 1593 30923
rect 1627 30920 1639 30923
rect 1762 30920 1768 30932
rect 1627 30892 1768 30920
rect 1627 30889 1639 30892
rect 1581 30883 1639 30889
rect 1762 30880 1768 30892
rect 1820 30880 1826 30932
rect 2133 30923 2191 30929
rect 2133 30889 2145 30923
rect 2179 30920 2191 30923
rect 2406 30920 2412 30932
rect 2179 30892 2412 30920
rect 2179 30889 2191 30892
rect 2133 30883 2191 30889
rect 2406 30880 2412 30892
rect 2464 30880 2470 30932
rect 2777 30923 2835 30929
rect 2777 30889 2789 30923
rect 2823 30920 2835 30923
rect 2958 30920 2964 30932
rect 2823 30892 2964 30920
rect 2823 30889 2835 30892
rect 2777 30883 2835 30889
rect 2958 30880 2964 30892
rect 3016 30880 3022 30932
rect 4706 30880 4712 30932
rect 4764 30920 4770 30932
rect 5442 30920 5448 30932
rect 4764 30892 5448 30920
rect 4764 30880 4770 30892
rect 5442 30880 5448 30892
rect 5500 30880 5506 30932
rect 934 30812 940 30864
rect 992 30852 998 30864
rect 992 30824 2360 30852
rect 992 30812 998 30824
rect 1486 30744 1492 30796
rect 1544 30784 1550 30796
rect 1946 30784 1952 30796
rect 1544 30756 1952 30784
rect 1544 30744 1550 30756
rect 1946 30744 1952 30756
rect 2004 30744 2010 30796
rect 1394 30716 1400 30728
rect 1355 30688 1400 30716
rect 1394 30676 1400 30688
rect 1452 30676 1458 30728
rect 2130 30716 2136 30728
rect 2043 30688 2136 30716
rect 2130 30676 2136 30688
rect 2188 30676 2194 30728
rect 2332 30725 2360 30824
rect 2317 30719 2375 30725
rect 2317 30685 2329 30719
rect 2363 30685 2375 30719
rect 2317 30679 2375 30685
rect 2498 30676 2504 30728
rect 2556 30716 2562 30728
rect 2777 30719 2835 30725
rect 2777 30716 2789 30719
rect 2556 30688 2789 30716
rect 2556 30676 2562 30688
rect 2777 30685 2789 30688
rect 2823 30685 2835 30719
rect 2777 30679 2835 30685
rect 2961 30719 3019 30725
rect 2961 30685 2973 30719
rect 3007 30716 3019 30719
rect 4065 30719 4123 30725
rect 3007 30688 3924 30716
rect 3007 30685 3019 30688
rect 2961 30679 3019 30685
rect 2148 30648 2176 30676
rect 2516 30648 2544 30676
rect 2148 30620 2544 30648
rect 3896 30589 3924 30688
rect 4065 30685 4077 30719
rect 4111 30716 4123 30719
rect 9766 30716 9772 30728
rect 4111 30688 9772 30716
rect 4111 30685 4123 30688
rect 4065 30679 4123 30685
rect 9766 30676 9772 30688
rect 9824 30676 9830 30728
rect 10134 30716 10140 30728
rect 10095 30688 10140 30716
rect 10134 30676 10140 30688
rect 10192 30676 10198 30728
rect 3881 30583 3939 30589
rect 3881 30549 3893 30583
rect 3927 30580 3939 30583
rect 5442 30580 5448 30592
rect 3927 30552 5448 30580
rect 3927 30549 3939 30552
rect 3881 30543 3939 30549
rect 5442 30540 5448 30552
rect 5500 30540 5506 30592
rect 9950 30580 9956 30592
rect 9911 30552 9956 30580
rect 9950 30540 9956 30552
rect 10008 30540 10014 30592
rect 1104 30490 10856 30512
rect 1104 30438 4213 30490
rect 4265 30438 4277 30490
rect 4329 30438 4341 30490
rect 4393 30438 4405 30490
rect 4457 30438 4469 30490
rect 4521 30438 7477 30490
rect 7529 30438 7541 30490
rect 7593 30438 7605 30490
rect 7657 30438 7669 30490
rect 7721 30438 7733 30490
rect 7785 30438 10856 30490
rect 1104 30416 10856 30438
rect 1578 30336 1584 30388
rect 1636 30376 1642 30388
rect 7190 30376 7196 30388
rect 1636 30348 7196 30376
rect 1636 30336 1642 30348
rect 7190 30336 7196 30348
rect 7248 30336 7254 30388
rect 5166 30308 5172 30320
rect 2608 30280 5172 30308
rect 1302 30200 1308 30252
rect 1360 30240 1366 30252
rect 1397 30243 1455 30249
rect 1397 30240 1409 30243
rect 1360 30212 1409 30240
rect 1360 30200 1366 30212
rect 1397 30209 1409 30212
rect 1443 30209 1455 30243
rect 1397 30203 1455 30209
rect 2314 30200 2320 30252
rect 2372 30240 2378 30252
rect 2608 30249 2636 30280
rect 5166 30268 5172 30280
rect 5224 30268 5230 30320
rect 2593 30243 2651 30249
rect 2593 30240 2605 30243
rect 2372 30212 2605 30240
rect 2372 30200 2378 30212
rect 2593 30209 2605 30212
rect 2639 30209 2651 30243
rect 2593 30203 2651 30209
rect 4065 30243 4123 30249
rect 4065 30209 4077 30243
rect 4111 30240 4123 30243
rect 9858 30240 9864 30252
rect 4111 30212 9864 30240
rect 4111 30209 4123 30212
rect 4065 30203 4123 30209
rect 9858 30200 9864 30212
rect 9916 30200 9922 30252
rect 10134 30240 10140 30252
rect 10095 30212 10140 30240
rect 10134 30200 10140 30212
rect 10192 30200 10198 30252
rect 2869 30175 2927 30181
rect 2869 30141 2881 30175
rect 2915 30172 2927 30175
rect 2958 30172 2964 30184
rect 2915 30144 2964 30172
rect 2915 30141 2927 30144
rect 2869 30135 2927 30141
rect 2958 30132 2964 30144
rect 3016 30132 3022 30184
rect 1581 30107 1639 30113
rect 1581 30073 1593 30107
rect 1627 30104 1639 30107
rect 1670 30104 1676 30116
rect 1627 30076 1676 30104
rect 1627 30073 1639 30076
rect 1581 30067 1639 30073
rect 1670 30064 1676 30076
rect 1728 30064 1734 30116
rect 3142 29996 3148 30048
rect 3200 30036 3206 30048
rect 3973 30039 4031 30045
rect 3973 30036 3985 30039
rect 3200 30008 3985 30036
rect 3200 29996 3206 30008
rect 3973 30005 3985 30008
rect 4019 30036 4031 30039
rect 5166 30036 5172 30048
rect 4019 30008 5172 30036
rect 4019 30005 4031 30008
rect 3973 29999 4031 30005
rect 5166 29996 5172 30008
rect 5224 29996 5230 30048
rect 9858 29996 9864 30048
rect 9916 30036 9922 30048
rect 9953 30039 10011 30045
rect 9953 30036 9965 30039
rect 9916 30008 9965 30036
rect 9916 29996 9922 30008
rect 9953 30005 9965 30008
rect 9999 30005 10011 30039
rect 9953 29999 10011 30005
rect 1104 29946 10856 29968
rect 1104 29894 2582 29946
rect 2634 29894 2646 29946
rect 2698 29894 2710 29946
rect 2762 29894 2774 29946
rect 2826 29894 2838 29946
rect 2890 29894 5845 29946
rect 5897 29894 5909 29946
rect 5961 29894 5973 29946
rect 6025 29894 6037 29946
rect 6089 29894 6101 29946
rect 6153 29894 9109 29946
rect 9161 29894 9173 29946
rect 9225 29894 9237 29946
rect 9289 29894 9301 29946
rect 9353 29894 9365 29946
rect 9417 29894 10856 29946
rect 1104 29872 10856 29894
rect 1578 29832 1584 29844
rect 1539 29804 1584 29832
rect 1578 29792 1584 29804
rect 1636 29792 1642 29844
rect 1762 29792 1768 29844
rect 1820 29832 1826 29844
rect 8478 29832 8484 29844
rect 1820 29804 8484 29832
rect 1820 29792 1826 29804
rect 8478 29792 8484 29804
rect 8536 29792 8542 29844
rect 2314 29696 2320 29708
rect 2275 29668 2320 29696
rect 2314 29656 2320 29668
rect 2372 29656 2378 29708
rect 2498 29656 2504 29708
rect 2556 29696 2562 29708
rect 2593 29699 2651 29705
rect 2593 29696 2605 29699
rect 2556 29668 2605 29696
rect 2556 29656 2562 29668
rect 2593 29665 2605 29668
rect 2639 29665 2651 29699
rect 2593 29659 2651 29665
rect 1394 29628 1400 29640
rect 1355 29600 1400 29628
rect 1394 29588 1400 29600
rect 1452 29588 1458 29640
rect 10134 29628 10140 29640
rect 10095 29600 10140 29628
rect 10134 29588 10140 29600
rect 10192 29588 10198 29640
rect 1670 29452 1676 29504
rect 1728 29492 1734 29504
rect 8294 29492 8300 29504
rect 1728 29464 8300 29492
rect 1728 29452 1734 29464
rect 8294 29452 8300 29464
rect 8352 29452 8358 29504
rect 9674 29452 9680 29504
rect 9732 29492 9738 29504
rect 9953 29495 10011 29501
rect 9953 29492 9965 29495
rect 9732 29464 9965 29492
rect 9732 29452 9738 29464
rect 9953 29461 9965 29464
rect 9999 29461 10011 29495
rect 9953 29455 10011 29461
rect 1104 29402 10856 29424
rect 1104 29350 4213 29402
rect 4265 29350 4277 29402
rect 4329 29350 4341 29402
rect 4393 29350 4405 29402
rect 4457 29350 4469 29402
rect 4521 29350 7477 29402
rect 7529 29350 7541 29402
rect 7593 29350 7605 29402
rect 7657 29350 7669 29402
rect 7721 29350 7733 29402
rect 7785 29350 10856 29402
rect 1104 29328 10856 29350
rect 1581 29291 1639 29297
rect 1581 29257 1593 29291
rect 1627 29288 1639 29291
rect 1670 29288 1676 29300
rect 1627 29260 1676 29288
rect 1627 29257 1639 29260
rect 1581 29251 1639 29257
rect 1670 29248 1676 29260
rect 1728 29248 1734 29300
rect 1854 29248 1860 29300
rect 1912 29288 1918 29300
rect 2225 29291 2283 29297
rect 2225 29288 2237 29291
rect 1912 29260 2237 29288
rect 1912 29248 1918 29260
rect 2225 29257 2237 29260
rect 2271 29257 2283 29291
rect 2225 29251 2283 29257
rect 2958 29220 2964 29232
rect 2148 29192 2964 29220
rect 1302 29112 1308 29164
rect 1360 29152 1366 29164
rect 2148 29161 2176 29192
rect 2958 29180 2964 29192
rect 3016 29180 3022 29232
rect 9674 29220 9680 29232
rect 9508 29192 9680 29220
rect 9508 29161 9536 29192
rect 9674 29180 9680 29192
rect 9732 29180 9738 29232
rect 1397 29155 1455 29161
rect 1397 29152 1409 29155
rect 1360 29124 1409 29152
rect 1360 29112 1366 29124
rect 1397 29121 1409 29124
rect 1443 29121 1455 29155
rect 1397 29115 1455 29121
rect 2133 29155 2191 29161
rect 2133 29121 2145 29155
rect 2179 29121 2191 29155
rect 2133 29115 2191 29121
rect 2317 29155 2375 29161
rect 2317 29121 2329 29155
rect 2363 29121 2375 29155
rect 2317 29115 2375 29121
rect 9493 29155 9551 29161
rect 9493 29121 9505 29155
rect 9539 29121 9551 29155
rect 9493 29115 9551 29121
rect 9585 29155 9643 29161
rect 9585 29121 9597 29155
rect 9631 29121 9643 29155
rect 9950 29152 9956 29164
rect 9911 29124 9956 29152
rect 9585 29115 9643 29121
rect 1210 29044 1216 29096
rect 1268 29084 1274 29096
rect 2332 29084 2360 29115
rect 1268 29056 2360 29084
rect 1268 29044 1274 29056
rect 3418 29044 3424 29096
rect 3476 29044 3482 29096
rect 3436 29016 3464 29044
rect 3344 28988 3464 29016
rect 9600 29016 9628 29115
rect 9950 29112 9956 29124
rect 10008 29112 10014 29164
rect 9950 29016 9956 29028
rect 9600 28988 9956 29016
rect 842 28908 848 28960
rect 900 28948 906 28960
rect 1486 28948 1492 28960
rect 900 28920 1492 28948
rect 900 28908 906 28920
rect 1486 28908 1492 28920
rect 1544 28908 1550 28960
rect 2038 28908 2044 28960
rect 2096 28948 2102 28960
rect 3344 28948 3372 28988
rect 9950 28976 9956 28988
rect 10008 28976 10014 29028
rect 2096 28920 3372 28948
rect 2096 28908 2102 28920
rect 3418 28908 3424 28960
rect 3476 28948 3482 28960
rect 4706 28948 4712 28960
rect 3476 28920 4712 28948
rect 3476 28908 3482 28920
rect 4706 28908 4712 28920
rect 4764 28908 4770 28960
rect 9858 28948 9864 28960
rect 9819 28920 9864 28948
rect 9858 28908 9864 28920
rect 9916 28908 9922 28960
rect 10137 28951 10195 28957
rect 10137 28917 10149 28951
rect 10183 28948 10195 28951
rect 10965 28951 11023 28957
rect 10965 28948 10977 28951
rect 10183 28920 10977 28948
rect 10183 28917 10195 28920
rect 10137 28911 10195 28917
rect 10965 28917 10977 28920
rect 11011 28917 11023 28951
rect 10965 28911 11023 28917
rect 1104 28858 10856 28880
rect 1104 28806 2582 28858
rect 2634 28806 2646 28858
rect 2698 28806 2710 28858
rect 2762 28806 2774 28858
rect 2826 28806 2838 28858
rect 2890 28806 5845 28858
rect 5897 28806 5909 28858
rect 5961 28806 5973 28858
rect 6025 28806 6037 28858
rect 6089 28806 6101 28858
rect 6153 28806 9109 28858
rect 9161 28806 9173 28858
rect 9225 28806 9237 28858
rect 9289 28806 9301 28858
rect 9353 28806 9365 28858
rect 9417 28806 10856 28858
rect 1104 28784 10856 28806
rect 1946 28704 1952 28756
rect 2004 28744 2010 28756
rect 2133 28747 2191 28753
rect 2133 28744 2145 28747
rect 2004 28716 2145 28744
rect 2004 28704 2010 28716
rect 2133 28713 2145 28716
rect 2179 28713 2191 28747
rect 2133 28707 2191 28713
rect 2777 28747 2835 28753
rect 2777 28713 2789 28747
rect 2823 28744 2835 28747
rect 3878 28744 3884 28756
rect 2823 28716 3884 28744
rect 2823 28713 2835 28716
rect 2777 28707 2835 28713
rect 3878 28704 3884 28716
rect 3936 28704 3942 28756
rect 9950 28744 9956 28756
rect 9911 28716 9956 28744
rect 9950 28704 9956 28716
rect 10008 28704 10014 28756
rect 1581 28679 1639 28685
rect 1581 28645 1593 28679
rect 1627 28676 1639 28679
rect 7006 28676 7012 28688
rect 1627 28648 7012 28676
rect 1627 28645 1639 28648
rect 1581 28639 1639 28645
rect 7006 28636 7012 28648
rect 7064 28636 7070 28688
rect 2148 28580 2820 28608
rect 1394 28540 1400 28552
rect 1355 28512 1400 28540
rect 1394 28500 1400 28512
rect 1452 28500 1458 28552
rect 2148 28549 2176 28580
rect 2792 28549 2820 28580
rect 2139 28543 2197 28549
rect 2139 28509 2151 28543
rect 2185 28509 2197 28543
rect 2139 28503 2197 28509
rect 2317 28543 2375 28549
rect 2317 28509 2329 28543
rect 2363 28509 2375 28543
rect 2317 28503 2375 28509
rect 2777 28543 2835 28549
rect 2777 28509 2789 28543
rect 2823 28540 2835 28543
rect 2866 28540 2872 28552
rect 2823 28512 2872 28540
rect 2823 28509 2835 28512
rect 2777 28503 2835 28509
rect 1026 28364 1032 28416
rect 1084 28404 1090 28416
rect 2332 28404 2360 28503
rect 2866 28500 2872 28512
rect 2924 28500 2930 28552
rect 2961 28543 3019 28549
rect 2961 28509 2973 28543
rect 3007 28540 3019 28543
rect 4706 28540 4712 28552
rect 3007 28512 4712 28540
rect 3007 28509 3019 28512
rect 2961 28503 3019 28509
rect 4706 28500 4712 28512
rect 4764 28500 4770 28552
rect 10134 28540 10140 28552
rect 10095 28512 10140 28540
rect 10134 28500 10140 28512
rect 10192 28500 10198 28552
rect 1084 28376 2360 28404
rect 1084 28364 1090 28376
rect 2498 28364 2504 28416
rect 2556 28404 2562 28416
rect 8754 28404 8760 28416
rect 2556 28376 8760 28404
rect 2556 28364 2562 28376
rect 8754 28364 8760 28376
rect 8812 28364 8818 28416
rect 1104 28314 10856 28336
rect 1104 28262 4213 28314
rect 4265 28262 4277 28314
rect 4329 28262 4341 28314
rect 4393 28262 4405 28314
rect 4457 28262 4469 28314
rect 4521 28262 7477 28314
rect 7529 28262 7541 28314
rect 7593 28262 7605 28314
rect 7657 28262 7669 28314
rect 7721 28262 7733 28314
rect 7785 28262 10856 28314
rect 1104 28240 10856 28262
rect 1581 28203 1639 28209
rect 1581 28169 1593 28203
rect 1627 28200 1639 28203
rect 1762 28200 1768 28212
rect 1627 28172 1768 28200
rect 1627 28169 1639 28172
rect 1581 28163 1639 28169
rect 1762 28160 1768 28172
rect 1820 28160 1826 28212
rect 2869 28203 2927 28209
rect 2869 28169 2881 28203
rect 2915 28200 2927 28203
rect 3510 28200 3516 28212
rect 2915 28172 3516 28200
rect 2915 28169 2927 28172
rect 2869 28163 2927 28169
rect 3510 28160 3516 28172
rect 3568 28160 3574 28212
rect 3878 28160 3884 28212
rect 3936 28200 3942 28212
rect 5074 28200 5080 28212
rect 3936 28172 5080 28200
rect 3936 28160 3942 28172
rect 5074 28160 5080 28172
rect 5132 28160 5138 28212
rect 934 28092 940 28144
rect 992 28132 998 28144
rect 1210 28132 1216 28144
rect 992 28104 1216 28132
rect 992 28092 998 28104
rect 1210 28092 1216 28104
rect 1268 28092 1274 28144
rect 2148 28104 2820 28132
rect 1302 28024 1308 28076
rect 1360 28064 1366 28076
rect 2148 28073 2176 28104
rect 2792 28073 2820 28104
rect 1397 28067 1455 28073
rect 1397 28064 1409 28067
rect 1360 28036 1409 28064
rect 1360 28024 1366 28036
rect 1397 28033 1409 28036
rect 1443 28033 1455 28067
rect 1397 28027 1455 28033
rect 2133 28067 2191 28073
rect 2133 28033 2145 28067
rect 2179 28033 2191 28067
rect 2133 28027 2191 28033
rect 2317 28067 2375 28073
rect 2317 28033 2329 28067
rect 2363 28033 2375 28067
rect 2317 28027 2375 28033
rect 2777 28067 2835 28073
rect 2777 28033 2789 28067
rect 2823 28064 2835 28067
rect 2866 28064 2872 28076
rect 2823 28036 2872 28064
rect 2823 28033 2835 28036
rect 2777 28027 2835 28033
rect 1210 27956 1216 28008
rect 1268 27996 1274 28008
rect 2332 27996 2360 28027
rect 2866 28024 2872 28036
rect 2924 28024 2930 28076
rect 2961 28067 3019 28073
rect 2961 28033 2973 28067
rect 3007 28064 3019 28067
rect 10134 28064 10140 28076
rect 3007 28036 4660 28064
rect 10095 28036 10140 28064
rect 3007 28033 3019 28036
rect 2961 28027 3019 28033
rect 4632 28008 4660 28036
rect 10134 28024 10140 28036
rect 10192 28024 10198 28076
rect 1268 27968 2360 27996
rect 1268 27956 1274 27968
rect 4614 27956 4620 28008
rect 4672 27956 4678 28008
rect 1578 27888 1584 27940
rect 1636 27928 1642 27940
rect 2133 27931 2191 27937
rect 2133 27928 2145 27931
rect 1636 27900 2145 27928
rect 1636 27888 1642 27900
rect 2133 27897 2145 27900
rect 2179 27897 2191 27931
rect 2133 27891 2191 27897
rect 9766 27820 9772 27872
rect 9824 27860 9830 27872
rect 9953 27863 10011 27869
rect 9953 27860 9965 27863
rect 9824 27832 9965 27860
rect 9824 27820 9830 27832
rect 9953 27829 9965 27832
rect 9999 27829 10011 27863
rect 9953 27823 10011 27829
rect 1104 27770 10856 27792
rect 1104 27718 2582 27770
rect 2634 27718 2646 27770
rect 2698 27718 2710 27770
rect 2762 27718 2774 27770
rect 2826 27718 2838 27770
rect 2890 27718 5845 27770
rect 5897 27718 5909 27770
rect 5961 27718 5973 27770
rect 6025 27718 6037 27770
rect 6089 27718 6101 27770
rect 6153 27718 9109 27770
rect 9161 27718 9173 27770
rect 9225 27718 9237 27770
rect 9289 27718 9301 27770
rect 9353 27718 9365 27770
rect 9417 27718 10856 27770
rect 1104 27696 10856 27718
rect 1857 27659 1915 27665
rect 1857 27625 1869 27659
rect 1903 27656 1915 27659
rect 2498 27656 2504 27668
rect 1903 27628 2504 27656
rect 1903 27625 1915 27628
rect 1857 27619 1915 27625
rect 2498 27616 2504 27628
rect 2556 27616 2562 27668
rect 2038 27548 2044 27600
rect 2096 27588 2102 27600
rect 3234 27588 3240 27600
rect 2096 27560 3240 27588
rect 2096 27548 2102 27560
rect 3234 27548 3240 27560
rect 3292 27548 3298 27600
rect 3418 27548 3424 27600
rect 3476 27588 3482 27600
rect 4522 27588 4528 27600
rect 3476 27560 4528 27588
rect 3476 27548 3482 27560
rect 4522 27548 4528 27560
rect 4580 27548 4586 27600
rect 658 27480 664 27532
rect 716 27520 722 27532
rect 2498 27520 2504 27532
rect 716 27492 2504 27520
rect 716 27480 722 27492
rect 2498 27480 2504 27492
rect 2556 27480 2562 27532
rect 106 27412 112 27464
rect 164 27452 170 27464
rect 2314 27452 2320 27464
rect 164 27424 2320 27452
rect 164 27412 170 27424
rect 2314 27412 2320 27424
rect 2372 27412 2378 27464
rect 10137 27455 10195 27461
rect 10137 27421 10149 27455
rect 10183 27452 10195 27455
rect 10226 27452 10232 27464
rect 10183 27424 10232 27452
rect 10183 27421 10195 27424
rect 10137 27415 10195 27421
rect 10226 27412 10232 27424
rect 10284 27412 10290 27464
rect 1946 27384 1952 27396
rect 1907 27356 1952 27384
rect 1946 27344 1952 27356
rect 2004 27344 2010 27396
rect 9858 27276 9864 27328
rect 9916 27316 9922 27328
rect 9953 27319 10011 27325
rect 9953 27316 9965 27319
rect 9916 27288 9965 27316
rect 9916 27276 9922 27288
rect 9953 27285 9965 27288
rect 9999 27285 10011 27319
rect 9953 27279 10011 27285
rect 1104 27226 10856 27248
rect 1104 27174 4213 27226
rect 4265 27174 4277 27226
rect 4329 27174 4341 27226
rect 4393 27174 4405 27226
rect 4457 27174 4469 27226
rect 4521 27174 7477 27226
rect 7529 27174 7541 27226
rect 7593 27174 7605 27226
rect 7657 27174 7669 27226
rect 7721 27174 7733 27226
rect 7785 27174 10856 27226
rect 1104 27152 10856 27174
rect 934 27004 940 27056
rect 992 27044 998 27056
rect 1210 27044 1216 27056
rect 992 27016 1216 27044
rect 992 27004 998 27016
rect 1210 27004 1216 27016
rect 1268 27004 1274 27056
rect 10042 26936 10048 26988
rect 10100 26976 10106 26988
rect 10137 26979 10195 26985
rect 10137 26976 10149 26979
rect 10100 26948 10149 26976
rect 10100 26936 10106 26948
rect 10137 26945 10149 26948
rect 10183 26945 10195 26979
rect 10137 26939 10195 26945
rect 9950 26772 9956 26784
rect 9911 26744 9956 26772
rect 9950 26732 9956 26744
rect 10008 26732 10014 26784
rect 1104 26682 10856 26704
rect 1104 26630 2582 26682
rect 2634 26630 2646 26682
rect 2698 26630 2710 26682
rect 2762 26630 2774 26682
rect 2826 26630 2838 26682
rect 2890 26630 5845 26682
rect 5897 26630 5909 26682
rect 5961 26630 5973 26682
rect 6025 26630 6037 26682
rect 6089 26630 6101 26682
rect 6153 26630 9109 26682
rect 9161 26630 9173 26682
rect 9225 26630 9237 26682
rect 9289 26630 9301 26682
rect 9353 26630 9365 26682
rect 9417 26630 10856 26682
rect 1104 26608 10856 26630
rect 1857 26571 1915 26577
rect 1857 26537 1869 26571
rect 1903 26568 1915 26571
rect 8662 26568 8668 26580
rect 1903 26540 8668 26568
rect 1903 26537 1915 26540
rect 1857 26531 1915 26537
rect 8662 26528 8668 26540
rect 8720 26528 8726 26580
rect 9858 26568 9864 26580
rect 9819 26540 9864 26568
rect 9858 26528 9864 26540
rect 9916 26528 9922 26580
rect 10045 26435 10103 26441
rect 10045 26401 10057 26435
rect 10091 26432 10103 26435
rect 10134 26432 10140 26444
rect 10091 26404 10140 26432
rect 10091 26401 10103 26404
rect 10045 26395 10103 26401
rect 10134 26392 10140 26404
rect 10192 26392 10198 26444
rect 9858 26364 9864 26376
rect 9819 26336 9864 26364
rect 9858 26324 9864 26336
rect 9916 26324 9922 26376
rect 1946 26296 1952 26308
rect 1907 26268 1952 26296
rect 1946 26256 1952 26268
rect 2004 26256 2010 26308
rect 10137 26299 10195 26305
rect 10137 26265 10149 26299
rect 10183 26296 10195 26299
rect 10965 26299 11023 26305
rect 10965 26296 10977 26299
rect 10183 26268 10977 26296
rect 10183 26265 10195 26268
rect 10137 26259 10195 26265
rect 10965 26265 10977 26268
rect 11011 26265 11023 26299
rect 10965 26259 11023 26265
rect 9677 26231 9735 26237
rect 9677 26197 9689 26231
rect 9723 26228 9735 26231
rect 10873 26231 10931 26237
rect 10873 26228 10885 26231
rect 9723 26200 10885 26228
rect 9723 26197 9735 26200
rect 9677 26191 9735 26197
rect 10873 26197 10885 26200
rect 10919 26197 10931 26231
rect 10873 26191 10931 26197
rect 1104 26138 10856 26160
rect 1104 26086 4213 26138
rect 4265 26086 4277 26138
rect 4329 26086 4341 26138
rect 4393 26086 4405 26138
rect 4457 26086 4469 26138
rect 4521 26086 7477 26138
rect 7529 26086 7541 26138
rect 7593 26086 7605 26138
rect 7657 26086 7669 26138
rect 7721 26086 7733 26138
rect 7785 26086 10856 26138
rect 1104 26064 10856 26086
rect 1857 26027 1915 26033
rect 1857 25993 1869 26027
rect 1903 26024 1915 26027
rect 8570 26024 8576 26036
rect 1903 25996 8576 26024
rect 1903 25993 1915 25996
rect 1857 25987 1915 25993
rect 8570 25984 8576 25996
rect 8628 25984 8634 26036
rect 10134 26024 10140 26036
rect 10095 25996 10140 26024
rect 10134 25984 10140 25996
rect 10192 25984 10198 26036
rect 9766 25956 9772 25968
rect 9727 25928 9772 25956
rect 9766 25916 9772 25928
rect 9824 25916 9830 25968
rect 9950 25956 9956 25968
rect 9911 25928 9956 25956
rect 9950 25916 9956 25928
rect 10008 25916 10014 25968
rect 1946 25888 1952 25900
rect 1907 25860 1952 25888
rect 1946 25848 1952 25860
rect 2004 25848 2010 25900
rect 1104 25594 10856 25616
rect 1104 25542 2582 25594
rect 2634 25542 2646 25594
rect 2698 25542 2710 25594
rect 2762 25542 2774 25594
rect 2826 25542 2838 25594
rect 2890 25542 5845 25594
rect 5897 25542 5909 25594
rect 5961 25542 5973 25594
rect 6025 25542 6037 25594
rect 6089 25542 6101 25594
rect 6153 25542 9109 25594
rect 9161 25542 9173 25594
rect 9225 25542 9237 25594
rect 9289 25542 9301 25594
rect 9353 25542 9365 25594
rect 9417 25542 10856 25594
rect 1104 25520 10856 25542
rect 1857 25483 1915 25489
rect 1857 25449 1869 25483
rect 1903 25480 1915 25483
rect 7282 25480 7288 25492
rect 1903 25452 7288 25480
rect 1903 25449 1915 25452
rect 1857 25443 1915 25449
rect 7282 25440 7288 25452
rect 7340 25440 7346 25492
rect 10134 25276 10140 25288
rect 10095 25248 10140 25276
rect 10134 25236 10140 25248
rect 10192 25236 10198 25288
rect 1946 25208 1952 25220
rect 1907 25180 1952 25208
rect 1946 25168 1952 25180
rect 2004 25168 2010 25220
rect 9766 25100 9772 25152
rect 9824 25140 9830 25152
rect 9953 25143 10011 25149
rect 9953 25140 9965 25143
rect 9824 25112 9965 25140
rect 9824 25100 9830 25112
rect 9953 25109 9965 25112
rect 9999 25109 10011 25143
rect 9953 25103 10011 25109
rect 1104 25050 10856 25072
rect 1104 24998 4213 25050
rect 4265 24998 4277 25050
rect 4329 24998 4341 25050
rect 4393 24998 4405 25050
rect 4457 24998 4469 25050
rect 4521 24998 7477 25050
rect 7529 24998 7541 25050
rect 7593 24998 7605 25050
rect 7657 24998 7669 25050
rect 7721 24998 7733 25050
rect 7785 24998 10856 25050
rect 1104 24976 10856 24998
rect 1946 24800 1952 24812
rect 1907 24772 1952 24800
rect 1946 24760 1952 24772
rect 2004 24760 2010 24812
rect 2501 24803 2559 24809
rect 2501 24769 2513 24803
rect 2547 24769 2559 24803
rect 2501 24763 2559 24769
rect 2516 24732 2544 24763
rect 2590 24760 2596 24812
rect 2648 24800 2654 24812
rect 2685 24803 2743 24809
rect 2685 24800 2697 24803
rect 2648 24772 2697 24800
rect 2648 24760 2654 24772
rect 2685 24769 2697 24772
rect 2731 24769 2743 24803
rect 2685 24763 2743 24769
rect 3145 24803 3203 24809
rect 3145 24769 3157 24803
rect 3191 24769 3203 24803
rect 3326 24800 3332 24812
rect 3287 24772 3332 24800
rect 3145 24763 3203 24769
rect 2958 24732 2964 24744
rect 2516 24704 2964 24732
rect 2958 24692 2964 24704
rect 3016 24732 3022 24744
rect 3160 24732 3188 24763
rect 3326 24760 3332 24772
rect 3384 24760 3390 24812
rect 10134 24800 10140 24812
rect 10095 24772 10140 24800
rect 10134 24760 10140 24772
rect 10192 24760 10198 24812
rect 3016 24704 3188 24732
rect 3016 24692 3022 24704
rect 1765 24667 1823 24673
rect 1765 24633 1777 24667
rect 1811 24664 1823 24667
rect 7098 24664 7104 24676
rect 1811 24636 7104 24664
rect 1811 24633 1823 24636
rect 1765 24627 1823 24633
rect 7098 24624 7104 24636
rect 7156 24624 7162 24676
rect 2498 24596 2504 24608
rect 2459 24568 2504 24596
rect 2498 24556 2504 24568
rect 2556 24556 2562 24608
rect 3145 24599 3203 24605
rect 3145 24565 3157 24599
rect 3191 24596 3203 24599
rect 3694 24596 3700 24608
rect 3191 24568 3700 24596
rect 3191 24565 3203 24568
rect 3145 24559 3203 24565
rect 3694 24556 3700 24568
rect 3752 24556 3758 24608
rect 9950 24596 9956 24608
rect 9911 24568 9956 24596
rect 9950 24556 9956 24568
rect 10008 24556 10014 24608
rect 1104 24506 10856 24528
rect 1104 24454 2582 24506
rect 2634 24454 2646 24506
rect 2698 24454 2710 24506
rect 2762 24454 2774 24506
rect 2826 24454 2838 24506
rect 2890 24454 5845 24506
rect 5897 24454 5909 24506
rect 5961 24454 5973 24506
rect 6025 24454 6037 24506
rect 6089 24454 6101 24506
rect 6153 24454 9109 24506
rect 9161 24454 9173 24506
rect 9225 24454 9237 24506
rect 9289 24454 9301 24506
rect 9353 24454 9365 24506
rect 9417 24454 10856 24506
rect 1104 24432 10856 24454
rect 1854 24392 1860 24404
rect 1815 24364 1860 24392
rect 1854 24352 1860 24364
rect 1912 24352 1918 24404
rect 2501 24191 2559 24197
rect 2501 24157 2513 24191
rect 2547 24157 2559 24191
rect 2501 24151 2559 24157
rect 2685 24191 2743 24197
rect 2685 24157 2697 24191
rect 2731 24188 2743 24191
rect 6270 24188 6276 24200
rect 2731 24160 6276 24188
rect 2731 24157 2743 24160
rect 2685 24151 2743 24157
rect 1946 24120 1952 24132
rect 1907 24092 1952 24120
rect 1946 24080 1952 24092
rect 2004 24080 2010 24132
rect 2516 24120 2544 24151
rect 6270 24148 6276 24160
rect 6328 24148 6334 24200
rect 10134 24188 10140 24200
rect 10095 24160 10140 24188
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 2866 24120 2872 24132
rect 2516 24092 2872 24120
rect 2866 24080 2872 24092
rect 2924 24080 2930 24132
rect 1762 24012 1768 24064
rect 1820 24052 1826 24064
rect 2593 24055 2651 24061
rect 2593 24052 2605 24055
rect 1820 24024 2605 24052
rect 1820 24012 1826 24024
rect 2593 24021 2605 24024
rect 2639 24021 2651 24055
rect 2593 24015 2651 24021
rect 9858 24012 9864 24064
rect 9916 24052 9922 24064
rect 9953 24055 10011 24061
rect 9953 24052 9965 24055
rect 9916 24024 9965 24052
rect 9916 24012 9922 24024
rect 9953 24021 9965 24024
rect 9999 24021 10011 24055
rect 9953 24015 10011 24021
rect 1104 23962 10856 23984
rect 1104 23910 4213 23962
rect 4265 23910 4277 23962
rect 4329 23910 4341 23962
rect 4393 23910 4405 23962
rect 4457 23910 4469 23962
rect 4521 23910 7477 23962
rect 7529 23910 7541 23962
rect 7593 23910 7605 23962
rect 7657 23910 7669 23962
rect 7721 23910 7733 23962
rect 7785 23910 10856 23962
rect 1104 23888 10856 23910
rect 2038 23780 2044 23792
rect 1999 23752 2044 23780
rect 2038 23740 2044 23752
rect 2096 23740 2102 23792
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 2777 23715 2835 23721
rect 2777 23681 2789 23715
rect 2823 23712 2835 23715
rect 2866 23712 2872 23724
rect 2823 23684 2872 23712
rect 2823 23681 2835 23684
rect 2777 23675 2835 23681
rect 2866 23672 2872 23684
rect 2924 23672 2930 23724
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3050 23712 3056 23724
rect 3007 23684 3056 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3050 23672 3056 23684
rect 3108 23672 3114 23724
rect 3421 23715 3479 23721
rect 3421 23681 3433 23715
rect 3467 23681 3479 23715
rect 3602 23712 3608 23724
rect 3563 23684 3608 23712
rect 3421 23675 3479 23681
rect 3436 23644 3464 23675
rect 3602 23672 3608 23684
rect 3660 23672 3666 23724
rect 9950 23712 9956 23724
rect 9911 23684 9956 23712
rect 9950 23672 9956 23684
rect 10008 23672 10014 23724
rect 3786 23644 3792 23656
rect 3436 23616 3792 23644
rect 3786 23604 3792 23616
rect 3844 23604 3850 23656
rect 2777 23579 2835 23585
rect 2777 23545 2789 23579
rect 2823 23576 2835 23579
rect 3326 23576 3332 23588
rect 2823 23548 3332 23576
rect 2823 23545 2835 23548
rect 2777 23539 2835 23545
rect 3326 23536 3332 23548
rect 3384 23536 3390 23588
rect 3142 23468 3148 23520
rect 3200 23508 3206 23520
rect 3421 23511 3479 23517
rect 3421 23508 3433 23511
rect 3200 23480 3433 23508
rect 3200 23468 3206 23480
rect 3421 23477 3433 23480
rect 3467 23477 3479 23511
rect 3421 23471 3479 23477
rect 10045 23511 10103 23517
rect 10045 23477 10057 23511
rect 10091 23508 10103 23511
rect 10134 23508 10140 23520
rect 10091 23480 10140 23508
rect 10091 23477 10103 23480
rect 10045 23471 10103 23477
rect 10134 23468 10140 23480
rect 10192 23468 10198 23520
rect 1104 23418 10856 23440
rect 1104 23366 2582 23418
rect 2634 23366 2646 23418
rect 2698 23366 2710 23418
rect 2762 23366 2774 23418
rect 2826 23366 2838 23418
rect 2890 23366 5845 23418
rect 5897 23366 5909 23418
rect 5961 23366 5973 23418
rect 6025 23366 6037 23418
rect 6089 23366 6101 23418
rect 6153 23366 9109 23418
rect 9161 23366 9173 23418
rect 9225 23366 9237 23418
rect 9289 23366 9301 23418
rect 9353 23366 9365 23418
rect 9417 23366 10856 23418
rect 1104 23344 10856 23366
rect 1857 23307 1915 23313
rect 1857 23273 1869 23307
rect 1903 23304 1915 23307
rect 7834 23304 7840 23316
rect 1903 23276 7840 23304
rect 1903 23273 1915 23276
rect 1857 23267 1915 23273
rect 7834 23264 7840 23276
rect 7892 23264 7898 23316
rect 9858 23304 9864 23316
rect 9819 23276 9864 23304
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 4890 23168 4896 23180
rect 2700 23140 4896 23168
rect 2700 23109 2728 23140
rect 4890 23128 4896 23140
rect 4948 23128 4954 23180
rect 9766 23168 9772 23180
rect 9727 23140 9772 23168
rect 9766 23128 9772 23140
rect 9824 23128 9830 23180
rect 9953 23171 10011 23177
rect 9953 23137 9965 23171
rect 9999 23168 10011 23171
rect 10042 23168 10048 23180
rect 9999 23140 10048 23168
rect 9999 23137 10011 23140
rect 9953 23131 10011 23137
rect 10042 23128 10048 23140
rect 10100 23128 10106 23180
rect 2501 23103 2559 23109
rect 2501 23069 2513 23103
rect 2547 23069 2559 23103
rect 2501 23063 2559 23069
rect 2685 23103 2743 23109
rect 2685 23069 2697 23103
rect 2731 23069 2743 23103
rect 3786 23100 3792 23112
rect 3747 23072 3792 23100
rect 2685 23063 2743 23069
rect 1946 23032 1952 23044
rect 1907 23004 1952 23032
rect 1946 22992 1952 23004
rect 2004 22992 2010 23044
rect 2516 23032 2544 23063
rect 3786 23060 3792 23072
rect 3844 23060 3850 23112
rect 3970 23100 3976 23112
rect 3931 23072 3976 23100
rect 3970 23060 3976 23072
rect 4028 23060 4034 23112
rect 9122 23100 9128 23112
rect 9083 23072 9128 23100
rect 9122 23060 9128 23072
rect 9180 23060 9186 23112
rect 2958 23032 2964 23044
rect 2516 23004 2964 23032
rect 2958 22992 2964 23004
rect 3016 22992 3022 23044
rect 10137 23035 10195 23041
rect 10137 23032 10149 23035
rect 9876 23004 10149 23032
rect 9876 22976 9904 23004
rect 10137 23001 10149 23004
rect 10183 23001 10195 23035
rect 10137 22995 10195 23001
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 2593 22967 2651 22973
rect 2593 22964 2605 22967
rect 1728 22936 2605 22964
rect 1728 22924 1734 22936
rect 2593 22933 2605 22936
rect 2639 22933 2651 22967
rect 2593 22927 2651 22933
rect 3050 22924 3056 22976
rect 3108 22964 3114 22976
rect 3881 22967 3939 22973
rect 3881 22964 3893 22967
rect 3108 22936 3893 22964
rect 3108 22924 3114 22936
rect 3881 22933 3893 22936
rect 3927 22933 3939 22967
rect 3881 22927 3939 22933
rect 9309 22967 9367 22973
rect 9309 22933 9321 22967
rect 9355 22964 9367 22967
rect 9582 22964 9588 22976
rect 9355 22936 9588 22964
rect 9355 22933 9367 22936
rect 9309 22927 9367 22933
rect 9582 22924 9588 22936
rect 9640 22924 9646 22976
rect 9858 22924 9864 22976
rect 9916 22924 9922 22976
rect 9950 22924 9956 22976
rect 10008 22964 10014 22976
rect 10045 22967 10103 22973
rect 10045 22964 10057 22967
rect 10008 22936 10057 22964
rect 10008 22924 10014 22936
rect 10045 22933 10057 22936
rect 10091 22933 10103 22967
rect 10045 22927 10103 22933
rect 1104 22874 10856 22896
rect 1104 22822 4213 22874
rect 4265 22822 4277 22874
rect 4329 22822 4341 22874
rect 4393 22822 4405 22874
rect 4457 22822 4469 22874
rect 4521 22822 7477 22874
rect 7529 22822 7541 22874
rect 7593 22822 7605 22874
rect 7657 22822 7669 22874
rect 7721 22822 7733 22874
rect 7785 22822 10856 22874
rect 1104 22800 10856 22822
rect 1857 22763 1915 22769
rect 1857 22729 1869 22763
rect 1903 22760 1915 22763
rect 7374 22760 7380 22772
rect 1903 22732 7380 22760
rect 1903 22729 1915 22732
rect 1857 22723 1915 22729
rect 7374 22720 7380 22732
rect 7432 22720 7438 22772
rect 9674 22760 9680 22772
rect 9635 22732 9680 22760
rect 9674 22720 9680 22732
rect 9732 22720 9738 22772
rect 1946 22624 1952 22636
rect 1907 22596 1952 22624
rect 1946 22584 1952 22596
rect 2004 22584 2010 22636
rect 2685 22627 2743 22633
rect 2685 22593 2697 22627
rect 2731 22624 2743 22627
rect 3234 22624 3240 22636
rect 2731 22596 3240 22624
rect 2731 22593 2743 22596
rect 2685 22587 2743 22593
rect 3234 22584 3240 22596
rect 3292 22584 3298 22636
rect 8846 22624 8852 22636
rect 8807 22596 8852 22624
rect 8846 22584 8852 22596
rect 8904 22584 8910 22636
rect 9950 22624 9956 22636
rect 9911 22596 9956 22624
rect 9950 22584 9956 22596
rect 10008 22584 10014 22636
rect 10134 22624 10140 22636
rect 10095 22596 10140 22624
rect 10134 22584 10140 22596
rect 10192 22584 10198 22636
rect 2958 22556 2964 22568
rect 2919 22528 2964 22556
rect 2958 22516 2964 22528
rect 3016 22516 3022 22568
rect 9585 22559 9643 22565
rect 9585 22525 9597 22559
rect 9631 22556 9643 22559
rect 10965 22559 11023 22565
rect 10965 22556 10977 22559
rect 9631 22528 10977 22556
rect 9631 22525 9643 22528
rect 9585 22519 9643 22525
rect 10965 22525 10977 22528
rect 11011 22525 11023 22559
rect 10965 22519 11023 22525
rect 9030 22420 9036 22432
rect 8991 22392 9036 22420
rect 9030 22380 9036 22392
rect 9088 22380 9094 22432
rect 1104 22330 10856 22352
rect 1104 22278 2582 22330
rect 2634 22278 2646 22330
rect 2698 22278 2710 22330
rect 2762 22278 2774 22330
rect 2826 22278 2838 22330
rect 2890 22278 5845 22330
rect 5897 22278 5909 22330
rect 5961 22278 5973 22330
rect 6025 22278 6037 22330
rect 6089 22278 6101 22330
rect 6153 22278 9109 22330
rect 9161 22278 9173 22330
rect 9225 22278 9237 22330
rect 9289 22278 9301 22330
rect 9353 22278 9365 22330
rect 9417 22278 10856 22330
rect 1104 22256 10856 22278
rect 10965 22151 11023 22157
rect 10965 22148 10977 22151
rect 10152 22120 10977 22148
rect 1765 22083 1823 22089
rect 1765 22049 1777 22083
rect 1811 22080 1823 22083
rect 8018 22080 8024 22092
rect 1811 22052 8024 22080
rect 1811 22049 1823 22052
rect 1765 22043 1823 22049
rect 8018 22040 8024 22052
rect 8076 22040 8082 22092
rect 9490 22080 9496 22092
rect 9451 22052 9496 22080
rect 9490 22040 9496 22052
rect 9548 22040 9554 22092
rect 1946 22012 1952 22024
rect 1907 21984 1952 22012
rect 1946 21972 1952 21984
rect 2004 21972 2010 22024
rect 2682 22021 2688 22024
rect 2507 22015 2565 22021
rect 2507 21981 2519 22015
rect 2553 21981 2565 22015
rect 2679 22012 2688 22021
rect 2643 21984 2688 22012
rect 2507 21975 2565 21981
rect 2679 21975 2688 21984
rect 2516 21944 2544 21975
rect 2682 21972 2688 21975
rect 2740 21972 2746 22024
rect 3602 21972 3608 22024
rect 3660 22012 3666 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3660 21984 3985 22012
rect 3660 21972 3666 21984
rect 3973 21981 3985 21984
rect 4019 22012 4031 22015
rect 9674 22012 9680 22024
rect 4019 21984 9680 22012
rect 4019 21981 4031 21984
rect 3973 21975 4031 21981
rect 9674 21972 9680 21984
rect 9732 21972 9738 22024
rect 9858 22012 9864 22024
rect 9819 21984 9864 22012
rect 9858 21972 9864 21984
rect 9916 21972 9922 22024
rect 10042 22012 10048 22024
rect 10003 21984 10048 22012
rect 10042 21972 10048 21984
rect 10100 21972 10106 22024
rect 10152 22021 10180 22120
rect 10965 22117 10977 22120
rect 11011 22117 11023 22151
rect 10965 22111 11023 22117
rect 10137 22015 10195 22021
rect 10137 21981 10149 22015
rect 10183 21981 10195 22015
rect 10137 21975 10195 21981
rect 2958 21944 2964 21956
rect 2516 21916 2964 21944
rect 2958 21904 2964 21916
rect 3016 21944 3022 21956
rect 3786 21944 3792 21956
rect 3016 21916 3792 21944
rect 3016 21904 3022 21916
rect 3786 21904 3792 21916
rect 3844 21904 3850 21956
rect 1946 21836 1952 21888
rect 2004 21876 2010 21888
rect 2593 21879 2651 21885
rect 2593 21876 2605 21879
rect 2004 21848 2605 21876
rect 2004 21836 2010 21848
rect 2593 21845 2605 21848
rect 2639 21845 2651 21879
rect 2593 21839 2651 21845
rect 3881 21879 3939 21885
rect 3881 21845 3893 21879
rect 3927 21876 3939 21879
rect 3970 21876 3976 21888
rect 3927 21848 3976 21876
rect 3927 21845 3939 21848
rect 3881 21839 3939 21845
rect 3970 21836 3976 21848
rect 4028 21836 4034 21888
rect 1104 21786 10856 21808
rect 1104 21734 4213 21786
rect 4265 21734 4277 21786
rect 4329 21734 4341 21786
rect 4393 21734 4405 21786
rect 4457 21734 4469 21786
rect 4521 21734 7477 21786
rect 7529 21734 7541 21786
rect 7593 21734 7605 21786
rect 7657 21734 7669 21786
rect 7721 21734 7733 21786
rect 7785 21734 10856 21786
rect 1104 21712 10856 21734
rect 566 21632 572 21684
rect 624 21672 630 21684
rect 3602 21672 3608 21684
rect 624 21644 3608 21672
rect 624 21632 630 21644
rect 3602 21632 3608 21644
rect 3660 21632 3666 21684
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 10137 21675 10195 21681
rect 10137 21672 10149 21675
rect 10100 21644 10149 21672
rect 10100 21632 10106 21644
rect 10137 21641 10149 21644
rect 10183 21641 10195 21675
rect 10137 21635 10195 21641
rect 1486 21564 1492 21616
rect 1544 21604 1550 21616
rect 2682 21604 2688 21616
rect 1544 21576 2688 21604
rect 1544 21564 1550 21576
rect 2682 21564 2688 21576
rect 2740 21564 2746 21616
rect 3237 21607 3295 21613
rect 3237 21573 3249 21607
rect 3283 21604 3295 21607
rect 3970 21604 3976 21616
rect 3283 21576 3976 21604
rect 3283 21573 3295 21576
rect 3237 21567 3295 21573
rect 3970 21564 3976 21576
rect 4028 21564 4034 21616
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 3142 21536 3148 21548
rect 1719 21508 3148 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 3142 21496 3148 21508
rect 3200 21496 3206 21548
rect 8938 21536 8944 21548
rect 8899 21508 8944 21536
rect 8938 21496 8944 21508
rect 8996 21496 9002 21548
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9766 21536 9772 21548
rect 9631 21508 9772 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9766 21496 9772 21508
rect 9824 21496 9830 21548
rect 9950 21536 9956 21548
rect 9911 21508 9956 21536
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 1486 21400 1492 21412
rect 1447 21372 1492 21400
rect 1486 21360 1492 21372
rect 1544 21360 1550 21412
rect 2958 21292 2964 21344
rect 3016 21332 3022 21344
rect 3142 21332 3148 21344
rect 3016 21304 3148 21332
rect 3016 21292 3022 21304
rect 3142 21292 3148 21304
rect 3200 21292 3206 21344
rect 3234 21292 3240 21344
rect 3292 21332 3298 21344
rect 3602 21332 3608 21344
rect 3292 21304 3608 21332
rect 3292 21292 3298 21304
rect 3602 21292 3608 21304
rect 3660 21332 3666 21344
rect 3881 21335 3939 21341
rect 3881 21332 3893 21335
rect 3660 21304 3893 21332
rect 3660 21292 3666 21304
rect 3881 21301 3893 21304
rect 3927 21301 3939 21335
rect 3881 21295 3939 21301
rect 9125 21335 9183 21341
rect 9125 21301 9137 21335
rect 9171 21332 9183 21335
rect 9582 21332 9588 21344
rect 9171 21304 9588 21332
rect 9171 21301 9183 21304
rect 9125 21295 9183 21301
rect 9582 21292 9588 21304
rect 9640 21292 9646 21344
rect 9858 21332 9864 21344
rect 9819 21304 9864 21332
rect 9858 21292 9864 21304
rect 9916 21292 9922 21344
rect 1104 21242 10856 21264
rect 1104 21190 2582 21242
rect 2634 21190 2646 21242
rect 2698 21190 2710 21242
rect 2762 21190 2774 21242
rect 2826 21190 2838 21242
rect 2890 21190 5845 21242
rect 5897 21190 5909 21242
rect 5961 21190 5973 21242
rect 6025 21190 6037 21242
rect 6089 21190 6101 21242
rect 6153 21190 9109 21242
rect 9161 21190 9173 21242
rect 9225 21190 9237 21242
rect 9289 21190 9301 21242
rect 9353 21190 9365 21242
rect 9417 21190 10856 21242
rect 1104 21168 10856 21190
rect 9217 21131 9275 21137
rect 9217 21097 9229 21131
rect 9263 21128 9275 21131
rect 9677 21131 9735 21137
rect 9677 21128 9689 21131
rect 9263 21100 9689 21128
rect 9263 21097 9275 21100
rect 9217 21091 9275 21097
rect 9677 21097 9689 21100
rect 9723 21097 9735 21131
rect 9677 21091 9735 21097
rect 9950 21088 9956 21140
rect 10008 21128 10014 21140
rect 10137 21131 10195 21137
rect 10137 21128 10149 21131
rect 10008 21100 10149 21128
rect 10008 21088 10014 21100
rect 10137 21097 10149 21100
rect 10183 21097 10195 21131
rect 10137 21091 10195 21097
rect 9582 20952 9588 21004
rect 9640 20992 9646 21004
rect 9769 20995 9827 21001
rect 9769 20992 9781 20995
rect 9640 20964 9781 20992
rect 9640 20952 9646 20964
rect 9769 20961 9781 20964
rect 9815 20961 9827 20995
rect 9769 20955 9827 20961
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 3050 20924 3056 20936
rect 1719 20896 3056 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 3050 20884 3056 20896
rect 3108 20884 3114 20936
rect 9030 20924 9036 20936
rect 8991 20896 9036 20924
rect 9030 20884 9036 20896
rect 9088 20884 9094 20936
rect 9674 20924 9680 20936
rect 9635 20896 9680 20924
rect 9674 20884 9680 20896
rect 9732 20884 9738 20936
rect 9953 20927 10011 20933
rect 9953 20893 9965 20927
rect 9999 20924 10011 20927
rect 10134 20924 10140 20936
rect 9999 20896 10140 20924
rect 9999 20893 10011 20896
rect 9953 20887 10011 20893
rect 10134 20884 10140 20896
rect 10192 20884 10198 20936
rect 750 20816 756 20868
rect 808 20856 814 20868
rect 2406 20856 2412 20868
rect 808 20828 2412 20856
rect 808 20816 814 20828
rect 2406 20816 2412 20828
rect 2464 20816 2470 20868
rect 1486 20788 1492 20800
rect 1447 20760 1492 20788
rect 1486 20748 1492 20760
rect 1544 20748 1550 20800
rect 1104 20698 10856 20720
rect 1104 20646 4213 20698
rect 4265 20646 4277 20698
rect 4329 20646 4341 20698
rect 4393 20646 4405 20698
rect 4457 20646 4469 20698
rect 4521 20646 7477 20698
rect 7529 20646 7541 20698
rect 7593 20646 7605 20698
rect 7657 20646 7669 20698
rect 7721 20646 7733 20698
rect 7785 20646 10856 20698
rect 1104 20624 10856 20646
rect 10042 20544 10048 20596
rect 10100 20584 10106 20596
rect 10137 20587 10195 20593
rect 10137 20584 10149 20587
rect 10100 20556 10149 20584
rect 10100 20544 10106 20556
rect 10137 20553 10149 20556
rect 10183 20553 10195 20587
rect 10137 20547 10195 20553
rect 9122 20476 9128 20528
rect 9180 20516 9186 20528
rect 9769 20519 9827 20525
rect 9769 20516 9781 20519
rect 9180 20488 9781 20516
rect 9180 20476 9186 20488
rect 9769 20485 9781 20488
rect 9815 20485 9827 20519
rect 9769 20479 9827 20485
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20448 1731 20451
rect 1946 20448 1952 20460
rect 1719 20420 1952 20448
rect 1719 20417 1731 20420
rect 1673 20411 1731 20417
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 9950 20448 9956 20460
rect 9911 20420 9956 20448
rect 9950 20408 9956 20420
rect 10008 20408 10014 20460
rect 1486 20312 1492 20324
rect 1447 20284 1492 20312
rect 1486 20272 1492 20284
rect 1544 20272 1550 20324
rect 1104 20154 10856 20176
rect 1104 20102 2582 20154
rect 2634 20102 2646 20154
rect 2698 20102 2710 20154
rect 2762 20102 2774 20154
rect 2826 20102 2838 20154
rect 2890 20102 5845 20154
rect 5897 20102 5909 20154
rect 5961 20102 5973 20154
rect 6025 20102 6037 20154
rect 6089 20102 6101 20154
rect 6153 20102 9109 20154
rect 9161 20102 9173 20154
rect 9225 20102 9237 20154
rect 9289 20102 9301 20154
rect 9353 20102 9365 20154
rect 9417 20102 10856 20154
rect 1104 20080 10856 20102
rect 9950 20040 9956 20052
rect 9911 20012 9956 20040
rect 9950 20000 9956 20012
rect 10008 20000 10014 20052
rect 1670 19836 1676 19848
rect 1631 19808 1676 19836
rect 1670 19796 1676 19808
rect 1728 19796 1734 19848
rect 10134 19836 10140 19848
rect 10095 19808 10140 19836
rect 10134 19796 10140 19808
rect 10192 19796 10198 19848
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 1104 19610 10856 19632
rect 1104 19558 4213 19610
rect 4265 19558 4277 19610
rect 4329 19558 4341 19610
rect 4393 19558 4405 19610
rect 4457 19558 4469 19610
rect 4521 19558 7477 19610
rect 7529 19558 7541 19610
rect 7593 19558 7605 19610
rect 7657 19558 7669 19610
rect 7721 19558 7733 19610
rect 7785 19558 10856 19610
rect 1104 19536 10856 19558
rect 9858 19456 9864 19508
rect 9916 19496 9922 19508
rect 9953 19499 10011 19505
rect 9953 19496 9965 19499
rect 9916 19468 9965 19496
rect 9916 19456 9922 19468
rect 9953 19465 9965 19468
rect 9999 19465 10011 19499
rect 9953 19459 10011 19465
rect 290 19388 296 19440
rect 348 19428 354 19440
rect 2038 19428 2044 19440
rect 348 19400 2044 19428
rect 348 19388 354 19400
rect 2038 19388 2044 19400
rect 2096 19388 2102 19440
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 3326 19360 3332 19372
rect 1719 19332 3332 19360
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 3326 19320 3332 19332
rect 3384 19320 3390 19372
rect 10137 19363 10195 19369
rect 10137 19329 10149 19363
rect 10183 19360 10195 19363
rect 10183 19332 10272 19360
rect 10183 19329 10195 19332
rect 10137 19323 10195 19329
rect 10244 19304 10272 19332
rect 10226 19252 10232 19304
rect 10284 19252 10290 19304
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 1104 19066 10856 19088
rect 1104 19014 2582 19066
rect 2634 19014 2646 19066
rect 2698 19014 2710 19066
rect 2762 19014 2774 19066
rect 2826 19014 2838 19066
rect 2890 19014 5845 19066
rect 5897 19014 5909 19066
rect 5961 19014 5973 19066
rect 6025 19014 6037 19066
rect 6089 19014 6101 19066
rect 6153 19014 9109 19066
rect 9161 19014 9173 19066
rect 9225 19014 9237 19066
rect 9289 19014 9301 19066
rect 9353 19014 9365 19066
rect 9417 19014 10856 19066
rect 1104 18992 10856 19014
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 1762 18748 1768 18760
rect 1719 18720 1768 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 1762 18708 1768 18720
rect 1820 18708 1826 18760
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 1104 18522 10856 18544
rect 1104 18470 4213 18522
rect 4265 18470 4277 18522
rect 4329 18470 4341 18522
rect 4393 18470 4405 18522
rect 4457 18470 4469 18522
rect 4521 18470 7477 18522
rect 7529 18470 7541 18522
rect 7593 18470 7605 18522
rect 7657 18470 7669 18522
rect 7721 18470 7733 18522
rect 7785 18470 10856 18522
rect 1104 18448 10856 18470
rect 3786 18340 3792 18352
rect 1688 18312 3792 18340
rect 1688 18281 1716 18312
rect 3786 18300 3792 18312
rect 3844 18300 3850 18352
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 1673 18235 1731 18241
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18241 2191 18275
rect 2314 18272 2320 18284
rect 2275 18244 2320 18272
rect 2133 18235 2191 18241
rect 2148 18204 2176 18235
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 2222 18204 2228 18216
rect 2148 18176 2228 18204
rect 2222 18164 2228 18176
rect 2280 18164 2286 18216
rect 382 18096 388 18148
rect 440 18136 446 18148
rect 2314 18136 2320 18148
rect 440 18108 2320 18136
rect 440 18096 446 18108
rect 2314 18096 2320 18108
rect 2372 18096 2378 18148
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 1670 18028 1676 18080
rect 1728 18068 1734 18080
rect 2133 18071 2191 18077
rect 2133 18068 2145 18071
rect 1728 18040 2145 18068
rect 1728 18028 1734 18040
rect 2133 18037 2145 18040
rect 2179 18037 2191 18071
rect 2133 18031 2191 18037
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 6730 18068 6736 18080
rect 3016 18040 6736 18068
rect 3016 18028 3022 18040
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 1104 17978 10856 18000
rect 1104 17926 2582 17978
rect 2634 17926 2646 17978
rect 2698 17926 2710 17978
rect 2762 17926 2774 17978
rect 2826 17926 2838 17978
rect 2890 17926 5845 17978
rect 5897 17926 5909 17978
rect 5961 17926 5973 17978
rect 6025 17926 6037 17978
rect 6089 17926 6101 17978
rect 6153 17926 9109 17978
rect 9161 17926 9173 17978
rect 9225 17926 9237 17978
rect 9289 17926 9301 17978
rect 9353 17926 9365 17978
rect 9417 17926 10856 17978
rect 1104 17904 10856 17926
rect 1946 17824 1952 17876
rect 2004 17864 2010 17876
rect 4062 17864 4068 17876
rect 2004 17836 4068 17864
rect 2004 17824 2010 17836
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 2498 17728 2504 17740
rect 1688 17700 2504 17728
rect 1688 17669 1716 17700
rect 2498 17688 2504 17700
rect 2556 17688 2562 17740
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17629 1731 17663
rect 1673 17623 1731 17629
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17660 2191 17663
rect 2222 17660 2228 17672
rect 2179 17632 2228 17660
rect 2179 17629 2191 17632
rect 2133 17623 2191 17629
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17660 2375 17663
rect 7926 17660 7932 17672
rect 2363 17632 7932 17660
rect 2363 17629 2375 17632
rect 2317 17623 2375 17629
rect 7926 17620 7932 17632
rect 7984 17620 7990 17672
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 1762 17484 1768 17536
rect 1820 17524 1826 17536
rect 2225 17527 2283 17533
rect 2225 17524 2237 17527
rect 1820 17496 2237 17524
rect 1820 17484 1826 17496
rect 2225 17493 2237 17496
rect 2271 17493 2283 17527
rect 2225 17487 2283 17493
rect 1104 17434 10856 17456
rect 1104 17382 4213 17434
rect 4265 17382 4277 17434
rect 4329 17382 4341 17434
rect 4393 17382 4405 17434
rect 4457 17382 4469 17434
rect 4521 17382 7477 17434
rect 7529 17382 7541 17434
rect 7593 17382 7605 17434
rect 7657 17382 7669 17434
rect 7721 17382 7733 17434
rect 7785 17382 10856 17434
rect 1104 17360 10856 17382
rect 3326 17280 3332 17332
rect 3384 17320 3390 17332
rect 5258 17320 5264 17332
rect 3384 17292 5264 17320
rect 3384 17280 3390 17292
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2222 17184 2228 17196
rect 2179 17156 2228 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 2222 17144 2228 17156
rect 2280 17144 2286 17196
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17184 2375 17187
rect 6362 17184 6368 17196
rect 2363 17156 6368 17184
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 2133 16983 2191 16989
rect 2133 16980 2145 16983
rect 1728 16952 2145 16980
rect 1728 16940 1734 16952
rect 2133 16949 2145 16952
rect 2179 16949 2191 16983
rect 2133 16943 2191 16949
rect 1104 16890 10856 16912
rect 1104 16838 2582 16890
rect 2634 16838 2646 16890
rect 2698 16838 2710 16890
rect 2762 16838 2774 16890
rect 2826 16838 2838 16890
rect 2890 16838 5845 16890
rect 5897 16838 5909 16890
rect 5961 16838 5973 16890
rect 6025 16838 6037 16890
rect 6089 16838 6101 16890
rect 6153 16838 9109 16890
rect 9161 16838 9173 16890
rect 9225 16838 9237 16890
rect 9289 16838 9301 16890
rect 9353 16838 9365 16890
rect 9417 16838 10856 16890
rect 1104 16816 10856 16838
rect 3786 16776 3792 16788
rect 2792 16748 3792 16776
rect 1854 16668 1860 16720
rect 1912 16708 1918 16720
rect 2133 16711 2191 16717
rect 2133 16708 2145 16711
rect 1912 16680 2145 16708
rect 1912 16668 1918 16680
rect 2133 16677 2145 16680
rect 2179 16677 2191 16711
rect 2133 16671 2191 16677
rect 2222 16640 2228 16652
rect 2135 16612 2228 16640
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 1762 16572 1768 16584
rect 1719 16544 1768 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 1762 16532 1768 16544
rect 1820 16532 1826 16584
rect 2148 16581 2176 16612
rect 2222 16600 2228 16612
rect 2280 16640 2286 16652
rect 2792 16640 2820 16748
rect 3786 16736 3792 16748
rect 3844 16736 3850 16788
rect 2958 16668 2964 16720
rect 3016 16668 3022 16720
rect 2280 16612 2820 16640
rect 2280 16600 2286 16612
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16541 2191 16575
rect 2133 16535 2191 16541
rect 2317 16575 2375 16581
rect 2317 16541 2329 16575
rect 2363 16572 2375 16575
rect 2406 16572 2412 16584
rect 2363 16544 2412 16572
rect 2363 16541 2375 16544
rect 2317 16535 2375 16541
rect 2406 16532 2412 16544
rect 2464 16532 2470 16584
rect 2792 16581 2820 16612
rect 2976 16581 3004 16668
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16541 2835 16575
rect 2777 16535 2835 16541
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16541 3019 16575
rect 2961 16535 3019 16541
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 2869 16439 2927 16445
rect 2869 16405 2881 16439
rect 2915 16436 2927 16439
rect 2958 16436 2964 16448
rect 2915 16408 2964 16436
rect 2915 16405 2927 16408
rect 2869 16399 2927 16405
rect 2958 16396 2964 16408
rect 3016 16396 3022 16448
rect 1104 16346 10856 16368
rect 1104 16294 4213 16346
rect 4265 16294 4277 16346
rect 4329 16294 4341 16346
rect 4393 16294 4405 16346
rect 4457 16294 4469 16346
rect 4521 16294 7477 16346
rect 7529 16294 7541 16346
rect 7593 16294 7605 16346
rect 7657 16294 7669 16346
rect 7721 16294 7733 16346
rect 7785 16294 10856 16346
rect 1104 16272 10856 16294
rect 6546 16164 6552 16176
rect 2332 16136 6552 16164
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 2332 16105 2360 16136
rect 6546 16124 6552 16136
rect 6604 16124 6610 16176
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16065 2191 16099
rect 2133 16059 2191 16065
rect 2317 16099 2375 16105
rect 2317 16065 2329 16099
rect 2363 16065 2375 16099
rect 2317 16059 2375 16065
rect 2777 16099 2835 16105
rect 2777 16065 2789 16099
rect 2823 16065 2835 16099
rect 2777 16059 2835 16065
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16096 3019 16099
rect 3694 16096 3700 16108
rect 3007 16068 3700 16096
rect 3007 16065 3019 16068
rect 2961 16059 3019 16065
rect 2148 16028 2176 16059
rect 2792 16028 2820 16059
rect 3694 16056 3700 16068
rect 3752 16056 3758 16108
rect 3234 16028 3240 16040
rect 2148 16000 3240 16028
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 1670 15852 1676 15904
rect 1728 15892 1734 15904
rect 2133 15895 2191 15901
rect 2133 15892 2145 15895
rect 1728 15864 2145 15892
rect 1728 15852 1734 15864
rect 2133 15861 2145 15864
rect 2179 15861 2191 15895
rect 2133 15855 2191 15861
rect 2777 15895 2835 15901
rect 2777 15861 2789 15895
rect 2823 15892 2835 15895
rect 3050 15892 3056 15904
rect 2823 15864 3056 15892
rect 2823 15861 2835 15864
rect 2777 15855 2835 15861
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 1104 15802 10856 15824
rect 1104 15750 2582 15802
rect 2634 15750 2646 15802
rect 2698 15750 2710 15802
rect 2762 15750 2774 15802
rect 2826 15750 2838 15802
rect 2890 15750 5845 15802
rect 5897 15750 5909 15802
rect 5961 15750 5973 15802
rect 6025 15750 6037 15802
rect 6089 15750 6101 15802
rect 6153 15750 9109 15802
rect 9161 15750 9173 15802
rect 9225 15750 9237 15802
rect 9289 15750 9301 15802
rect 9353 15750 9365 15802
rect 9417 15750 10856 15802
rect 1104 15728 10856 15750
rect 2958 15620 2964 15632
rect 1688 15592 2964 15620
rect 1688 15493 1716 15592
rect 2958 15580 2964 15592
rect 3016 15580 3022 15632
rect 2038 15512 2044 15564
rect 2096 15552 2102 15564
rect 3234 15552 3240 15564
rect 2096 15524 2360 15552
rect 2096 15512 2102 15524
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 2130 15484 2136 15496
rect 2091 15456 2136 15484
rect 1673 15447 1731 15453
rect 2130 15444 2136 15456
rect 2188 15444 2194 15496
rect 2332 15493 2360 15524
rect 2792 15524 3240 15552
rect 2792 15493 2820 15524
rect 3234 15512 3240 15524
rect 3292 15552 3298 15564
rect 3418 15552 3424 15564
rect 3292 15524 3424 15552
rect 3292 15512 3298 15524
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15453 2375 15487
rect 2317 15447 2375 15453
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15453 2835 15487
rect 2777 15447 2835 15453
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 6822 15484 6828 15496
rect 3007 15456 6828 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 6822 15444 6828 15456
rect 6880 15444 6886 15496
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 2222 15348 2228 15360
rect 2183 15320 2228 15348
rect 2222 15308 2228 15320
rect 2280 15308 2286 15360
rect 2869 15351 2927 15357
rect 2869 15317 2881 15351
rect 2915 15348 2927 15351
rect 3234 15348 3240 15360
rect 2915 15320 3240 15348
rect 2915 15317 2927 15320
rect 2869 15311 2927 15317
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 1104 15258 10856 15280
rect 1104 15206 4213 15258
rect 4265 15206 4277 15258
rect 4329 15206 4341 15258
rect 4393 15206 4405 15258
rect 4457 15206 4469 15258
rect 4521 15206 7477 15258
rect 7529 15206 7541 15258
rect 7593 15206 7605 15258
rect 7657 15206 7669 15258
rect 7721 15206 7733 15258
rect 7785 15206 10856 15258
rect 1104 15184 10856 15206
rect 2148 15048 2820 15076
rect 2148 15020 2176 15048
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 1854 15008 1860 15020
rect 1719 14980 1860 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 2792 15017 2820 15048
rect 3510 15036 3516 15088
rect 3568 15076 3574 15088
rect 3568 15048 3648 15076
rect 3568 15036 3574 15048
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 14977 2375 15011
rect 2317 14971 2375 14977
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 14977 2835 15011
rect 2777 14971 2835 14977
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 3326 15008 3332 15020
rect 3007 14980 3332 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 2332 14940 2360 14971
rect 3326 14968 3332 14980
rect 3384 14968 3390 15020
rect 3418 14968 3424 15020
rect 3476 15008 3482 15020
rect 3620 15017 3648 15048
rect 3605 15011 3663 15017
rect 3476 14980 3521 15008
rect 3476 14968 3482 14980
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 6178 14940 6184 14952
rect 2332 14912 6184 14940
rect 6178 14900 6184 14912
rect 6236 14900 6242 14952
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 2133 14807 2191 14813
rect 2133 14804 2145 14807
rect 1820 14776 2145 14804
rect 1820 14764 1826 14776
rect 2133 14773 2145 14776
rect 2179 14773 2191 14807
rect 2133 14767 2191 14773
rect 2777 14807 2835 14813
rect 2777 14773 2789 14807
rect 2823 14804 2835 14807
rect 3050 14804 3056 14816
rect 2823 14776 3056 14804
rect 2823 14773 2835 14776
rect 2777 14767 2835 14773
rect 3050 14764 3056 14776
rect 3108 14764 3114 14816
rect 3418 14804 3424 14816
rect 3379 14776 3424 14804
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 1104 14714 10856 14736
rect 1104 14662 2582 14714
rect 2634 14662 2646 14714
rect 2698 14662 2710 14714
rect 2762 14662 2774 14714
rect 2826 14662 2838 14714
rect 2890 14662 5845 14714
rect 5897 14662 5909 14714
rect 5961 14662 5973 14714
rect 6025 14662 6037 14714
rect 6089 14662 6101 14714
rect 6153 14662 9109 14714
rect 9161 14662 9173 14714
rect 9225 14662 9237 14714
rect 9289 14662 9301 14714
rect 9353 14662 9365 14714
rect 9417 14662 10856 14714
rect 1104 14640 10856 14662
rect 2958 14532 2964 14544
rect 1688 14504 2964 14532
rect 1688 14405 1716 14504
rect 2958 14492 2964 14504
rect 3016 14492 3022 14544
rect 5626 14464 5632 14476
rect 2976 14436 5632 14464
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 2130 14396 2136 14408
rect 2043 14368 2136 14396
rect 1673 14359 1731 14365
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 2314 14396 2320 14408
rect 2275 14368 2320 14396
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 2498 14356 2504 14408
rect 2556 14396 2562 14408
rect 2976 14405 3004 14436
rect 5626 14424 5632 14436
rect 5684 14424 5690 14476
rect 2777 14399 2835 14405
rect 2777 14396 2789 14399
rect 2556 14368 2789 14396
rect 2556 14356 2562 14368
rect 2777 14365 2789 14368
rect 2823 14365 2835 14399
rect 2777 14359 2835 14365
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14365 3019 14399
rect 2961 14359 3019 14365
rect 3326 14356 3332 14408
rect 3384 14396 3390 14408
rect 3789 14399 3847 14405
rect 3789 14396 3801 14399
rect 3384 14368 3801 14396
rect 3384 14356 3390 14368
rect 3789 14365 3801 14368
rect 3835 14365 3847 14399
rect 3789 14359 3847 14365
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 3936 14368 3985 14396
rect 3936 14356 3942 14368
rect 3973 14365 3985 14368
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 2148 14328 2176 14356
rect 2516 14328 2544 14356
rect 2148 14300 2544 14328
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2130 14220 2136 14272
rect 2188 14260 2194 14272
rect 2225 14263 2283 14269
rect 2225 14260 2237 14263
rect 2188 14232 2237 14260
rect 2188 14220 2194 14232
rect 2225 14229 2237 14232
rect 2271 14229 2283 14263
rect 2225 14223 2283 14229
rect 2869 14263 2927 14269
rect 2869 14229 2881 14263
rect 2915 14260 2927 14263
rect 2958 14260 2964 14272
rect 2915 14232 2964 14260
rect 2915 14229 2927 14232
rect 2869 14223 2927 14229
rect 2958 14220 2964 14232
rect 3016 14220 3022 14272
rect 3878 14260 3884 14272
rect 3839 14232 3884 14260
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 1104 14170 10856 14192
rect 1104 14118 4213 14170
rect 4265 14118 4277 14170
rect 4329 14118 4341 14170
rect 4393 14118 4405 14170
rect 4457 14118 4469 14170
rect 4521 14118 7477 14170
rect 7529 14118 7541 14170
rect 7593 14118 7605 14170
rect 7657 14118 7669 14170
rect 7721 14118 7733 14170
rect 7785 14118 10856 14170
rect 1104 14096 10856 14118
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 3878 13920 3884 13932
rect 1719 13892 3884 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 3878 13880 3884 13892
rect 3936 13880 3942 13932
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13852 3295 13855
rect 3326 13852 3332 13864
rect 3283 13824 3332 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 3513 13855 3571 13861
rect 3513 13821 3525 13855
rect 3559 13852 3571 13855
rect 3602 13852 3608 13864
rect 3559 13824 3608 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 474 13744 480 13796
rect 532 13784 538 13796
rect 1394 13784 1400 13796
rect 532 13756 1400 13784
rect 532 13744 538 13756
rect 1394 13744 1400 13756
rect 1452 13744 1458 13796
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 1104 13626 10856 13648
rect 1104 13574 2582 13626
rect 2634 13574 2646 13626
rect 2698 13574 2710 13626
rect 2762 13574 2774 13626
rect 2826 13574 2838 13626
rect 2890 13574 5845 13626
rect 5897 13574 5909 13626
rect 5961 13574 5973 13626
rect 6025 13574 6037 13626
rect 6089 13574 6101 13626
rect 6153 13574 9109 13626
rect 9161 13574 9173 13626
rect 9225 13574 9237 13626
rect 9289 13574 9301 13626
rect 9353 13574 9365 13626
rect 9417 13574 10856 13626
rect 1104 13552 10856 13574
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 2639 13515 2697 13521
rect 2639 13512 2651 13515
rect 2556 13484 2651 13512
rect 2556 13472 2562 13484
rect 2639 13481 2651 13484
rect 2685 13481 2697 13515
rect 2639 13475 2697 13481
rect 3418 13444 3424 13456
rect 1688 13416 3424 13444
rect 1688 13317 1716 13416
rect 3418 13404 3424 13416
rect 3476 13404 3482 13456
rect 2409 13379 2467 13385
rect 2409 13345 2421 13379
rect 2455 13376 2467 13379
rect 2455 13348 2774 13376
rect 2455 13345 2467 13348
rect 2409 13339 2467 13345
rect 2746 13320 2774 13348
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13277 1731 13311
rect 2746 13308 2780 13320
rect 2687 13280 2780 13308
rect 1673 13271 1731 13277
rect 2774 13268 2780 13280
rect 2832 13308 2838 13320
rect 3602 13308 3608 13320
rect 2832 13280 3608 13308
rect 2832 13268 2838 13280
rect 3602 13268 3608 13280
rect 3660 13268 3666 13320
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 1104 13082 10856 13104
rect 1104 13030 4213 13082
rect 4265 13030 4277 13082
rect 4329 13030 4341 13082
rect 4393 13030 4405 13082
rect 4457 13030 4469 13082
rect 4521 13030 7477 13082
rect 7529 13030 7541 13082
rect 7593 13030 7605 13082
rect 7657 13030 7669 13082
rect 7721 13030 7733 13082
rect 7785 13030 10856 13082
rect 1104 13008 10856 13030
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12832 2743 12835
rect 2774 12832 2780 12844
rect 2731 12804 2780 12832
rect 2731 12801 2743 12804
rect 2685 12795 2743 12801
rect 2774 12792 2780 12804
rect 2832 12792 2838 12844
rect 2961 12835 3019 12841
rect 2961 12801 2973 12835
rect 3007 12832 3019 12835
rect 3786 12832 3792 12844
rect 3007 12804 3792 12832
rect 3007 12801 3019 12804
rect 2961 12795 3019 12801
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 1118 12724 1124 12776
rect 1176 12764 1182 12776
rect 3326 12764 3332 12776
rect 1176 12736 3332 12764
rect 1176 12724 1182 12736
rect 3326 12724 3332 12736
rect 3384 12724 3390 12776
rect 1486 12628 1492 12640
rect 1447 12600 1492 12628
rect 1486 12588 1492 12600
rect 1544 12588 1550 12640
rect 3970 12588 3976 12640
rect 4028 12628 4034 12640
rect 5442 12628 5448 12640
rect 4028 12600 5448 12628
rect 4028 12588 4034 12600
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 1104 12538 10856 12560
rect 1104 12486 2582 12538
rect 2634 12486 2646 12538
rect 2698 12486 2710 12538
rect 2762 12486 2774 12538
rect 2826 12486 2838 12538
rect 2890 12486 5845 12538
rect 5897 12486 5909 12538
rect 5961 12486 5973 12538
rect 6025 12486 6037 12538
rect 6089 12486 6101 12538
rect 6153 12486 9109 12538
rect 9161 12486 9173 12538
rect 9225 12486 9237 12538
rect 9289 12486 9301 12538
rect 9353 12486 9365 12538
rect 9417 12486 10856 12538
rect 1104 12464 10856 12486
rect 198 12384 204 12436
rect 256 12424 262 12436
rect 1578 12424 1584 12436
rect 256 12396 1584 12424
rect 256 12384 262 12396
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 3234 12220 3240 12232
rect 1719 12192 3240 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 1104 11994 10856 12016
rect 1104 11942 4213 11994
rect 4265 11942 4277 11994
rect 4329 11942 4341 11994
rect 4393 11942 4405 11994
rect 4457 11942 4469 11994
rect 4521 11942 7477 11994
rect 7529 11942 7541 11994
rect 7593 11942 7605 11994
rect 7657 11942 7669 11994
rect 7721 11942 7733 11994
rect 7785 11942 10856 11994
rect 1104 11920 10856 11942
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 3050 11744 3056 11756
rect 1719 11716 3056 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 1486 11540 1492 11552
rect 1447 11512 1492 11540
rect 1486 11500 1492 11512
rect 1544 11500 1550 11552
rect 1104 11450 10856 11472
rect 1104 11398 2582 11450
rect 2634 11398 2646 11450
rect 2698 11398 2710 11450
rect 2762 11398 2774 11450
rect 2826 11398 2838 11450
rect 2890 11398 5845 11450
rect 5897 11398 5909 11450
rect 5961 11398 5973 11450
rect 6025 11398 6037 11450
rect 6089 11398 6101 11450
rect 6153 11398 9109 11450
rect 9161 11398 9173 11450
rect 9225 11398 9237 11450
rect 9289 11398 9301 11450
rect 9353 11398 9365 11450
rect 9417 11398 10856 11450
rect 1104 11376 10856 11398
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 2222 11132 2228 11144
rect 1719 11104 2228 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 2222 11092 2228 11104
rect 2280 11092 2286 11144
rect 3418 11024 3424 11076
rect 3476 11064 3482 11076
rect 5166 11064 5172 11076
rect 3476 11036 5172 11064
rect 3476 11024 3482 11036
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 1486 10996 1492 11008
rect 1447 10968 1492 10996
rect 1486 10956 1492 10968
rect 1544 10956 1550 11008
rect 1104 10906 10856 10928
rect 1104 10854 4213 10906
rect 4265 10854 4277 10906
rect 4329 10854 4341 10906
rect 4393 10854 4405 10906
rect 4457 10854 4469 10906
rect 4521 10854 7477 10906
rect 7529 10854 7541 10906
rect 7593 10854 7605 10906
rect 7657 10854 7669 10906
rect 7721 10854 7733 10906
rect 7785 10854 10856 10906
rect 1104 10832 10856 10854
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2958 10656 2964 10668
rect 1719 10628 2964 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 1104 10362 10856 10384
rect 1104 10310 2582 10362
rect 2634 10310 2646 10362
rect 2698 10310 2710 10362
rect 2762 10310 2774 10362
rect 2826 10310 2838 10362
rect 2890 10310 5845 10362
rect 5897 10310 5909 10362
rect 5961 10310 5973 10362
rect 6025 10310 6037 10362
rect 6089 10310 6101 10362
rect 6153 10310 9109 10362
rect 9161 10310 9173 10362
rect 9225 10310 9237 10362
rect 9289 10310 9301 10362
rect 9353 10310 9365 10362
rect 9417 10310 10856 10362
rect 1104 10288 10856 10310
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 3602 10112 3608 10124
rect 3283 10084 3608 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 3602 10072 3608 10084
rect 3660 10072 3666 10124
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 1762 10044 1768 10056
rect 1719 10016 1768 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3050 10044 3056 10056
rect 3007 10016 3056 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 1486 9908 1492 9920
rect 1447 9880 1492 9908
rect 1486 9868 1492 9880
rect 1544 9868 1550 9920
rect 1104 9818 10856 9840
rect 1104 9766 4213 9818
rect 4265 9766 4277 9818
rect 4329 9766 4341 9818
rect 4393 9766 4405 9818
rect 4457 9766 4469 9818
rect 4521 9766 7477 9818
rect 7529 9766 7541 9818
rect 7593 9766 7605 9818
rect 7657 9766 7669 9818
rect 7721 9766 7733 9818
rect 7785 9766 10856 9818
rect 1104 9744 10856 9766
rect 1670 9568 1676 9580
rect 1631 9540 1676 9568
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 1486 9364 1492 9376
rect 1447 9336 1492 9364
rect 1486 9324 1492 9336
rect 1544 9324 1550 9376
rect 2314 9364 2320 9376
rect 2275 9336 2320 9364
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 1104 9274 10856 9296
rect 1104 9222 2582 9274
rect 2634 9222 2646 9274
rect 2698 9222 2710 9274
rect 2762 9222 2774 9274
rect 2826 9222 2838 9274
rect 2890 9222 5845 9274
rect 5897 9222 5909 9274
rect 5961 9222 5973 9274
rect 6025 9222 6037 9274
rect 6089 9222 6101 9274
rect 6153 9222 9109 9274
rect 9161 9222 9173 9274
rect 9225 9222 9237 9274
rect 9289 9222 9301 9274
rect 9353 9222 9365 9274
rect 9417 9222 10856 9274
rect 1104 9200 10856 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 1728 9132 2973 9160
rect 1728 9120 1734 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 2961 9123 3019 9129
rect 934 9052 940 9104
rect 992 9092 998 9104
rect 2314 9092 2320 9104
rect 992 9064 2320 9092
rect 992 9052 998 9064
rect 2314 9052 2320 9064
rect 2372 9052 2378 9104
rect 1394 8984 1400 9036
rect 1452 9024 1458 9036
rect 1452 8996 2360 9024
rect 1452 8984 1458 8996
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 2222 8956 2228 8968
rect 1719 8928 2228 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 2332 8965 2360 8996
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2961 8959 3019 8965
rect 2961 8956 2973 8959
rect 2547 8928 2973 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2961 8925 2973 8928
rect 3007 8956 3019 8959
rect 3050 8956 3056 8968
rect 3007 8928 3056 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8956 3203 8959
rect 3326 8956 3332 8968
rect 3191 8928 3332 8956
rect 3191 8925 3203 8928
rect 3145 8919 3203 8925
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 1394 8780 1400 8832
rect 1452 8820 1458 8832
rect 1489 8823 1547 8829
rect 1489 8820 1501 8823
rect 1452 8792 1501 8820
rect 1452 8780 1458 8792
rect 1489 8789 1501 8792
rect 1535 8789 1547 8823
rect 1489 8783 1547 8789
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 2409 8823 2467 8829
rect 2409 8820 2421 8823
rect 1728 8792 2421 8820
rect 1728 8780 1734 8792
rect 2409 8789 2421 8792
rect 2455 8789 2467 8823
rect 2409 8783 2467 8789
rect 1104 8730 10856 8752
rect 1104 8678 4213 8730
rect 4265 8678 4277 8730
rect 4329 8678 4341 8730
rect 4393 8678 4405 8730
rect 4457 8678 4469 8730
rect 4521 8678 7477 8730
rect 7529 8678 7541 8730
rect 7593 8678 7605 8730
rect 7657 8678 7669 8730
rect 7721 8678 7733 8730
rect 7785 8678 10856 8730
rect 1104 8656 10856 8678
rect 2222 8576 2228 8628
rect 2280 8616 2286 8628
rect 3513 8619 3571 8625
rect 3513 8616 3525 8619
rect 2280 8588 3525 8616
rect 2280 8576 2286 8588
rect 3513 8585 3525 8588
rect 3559 8585 3571 8619
rect 3513 8579 3571 8585
rect 1578 8508 1584 8560
rect 1636 8548 1642 8560
rect 3050 8548 3056 8560
rect 1636 8520 2360 8548
rect 1636 8508 1642 8520
rect 1670 8480 1676 8492
rect 1631 8452 1676 8480
rect 1670 8440 1676 8452
rect 1728 8440 1734 8492
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 2332 8489 2360 8520
rect 2792 8520 3056 8548
rect 2792 8489 2820 8520
rect 3050 8508 3056 8520
rect 3108 8548 3114 8560
rect 3108 8520 3464 8548
rect 3108 8508 3114 8520
rect 3436 8489 3464 8520
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8449 2835 8483
rect 2777 8443 2835 8449
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8480 3479 8483
rect 3510 8480 3516 8492
rect 3467 8452 3516 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 2976 8412 3004 8443
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 4982 8480 4988 8492
rect 3651 8452 4988 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5350 8412 5356 8424
rect 2976 8384 5356 8412
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 1670 8304 1676 8356
rect 1728 8344 1734 8356
rect 2133 8347 2191 8353
rect 2133 8344 2145 8347
rect 1728 8316 2145 8344
rect 1728 8304 1734 8316
rect 2133 8313 2145 8316
rect 2179 8313 2191 8347
rect 2133 8307 2191 8313
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8276 2835 8279
rect 2958 8276 2964 8288
rect 2823 8248 2964 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 1104 8186 10856 8208
rect 1104 8134 2582 8186
rect 2634 8134 2646 8186
rect 2698 8134 2710 8186
rect 2762 8134 2774 8186
rect 2826 8134 2838 8186
rect 2890 8134 5845 8186
rect 5897 8134 5909 8186
rect 5961 8134 5973 8186
rect 6025 8134 6037 8186
rect 6089 8134 6101 8186
rect 6153 8134 9109 8186
rect 9161 8134 9173 8186
rect 9225 8134 9237 8186
rect 9289 8134 9301 8186
rect 9353 8134 9365 8186
rect 9417 8134 10856 8186
rect 1104 8112 10856 8134
rect 2958 8004 2964 8016
rect 2746 7976 2964 8004
rect 2746 7936 2774 7976
rect 2958 7964 2964 7976
rect 3016 7964 3022 8016
rect 5534 7936 5540 7948
rect 1688 7908 2774 7936
rect 2976 7908 5540 7936
rect 1688 7877 1716 7908
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 2130 7868 2136 7880
rect 2043 7840 2136 7868
rect 1673 7831 1731 7837
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 2314 7868 2320 7880
rect 2275 7840 2320 7868
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 2976 7877 3004 7908
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2961 7871 3019 7877
rect 2823 7840 2857 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 2148 7800 2176 7828
rect 2792 7800 2820 7831
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3568 7840 3801 7868
rect 3568 7828 3574 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4798 7868 4804 7880
rect 4019 7840 4804 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 3234 7800 3240 7812
rect 2148 7772 3240 7800
rect 3234 7760 3240 7772
rect 3292 7760 3298 7812
rect 1302 7692 1308 7744
rect 1360 7732 1366 7744
rect 1489 7735 1547 7741
rect 1489 7732 1501 7735
rect 1360 7704 1501 7732
rect 1360 7692 1366 7704
rect 1489 7701 1501 7704
rect 1535 7701 1547 7735
rect 2222 7732 2228 7744
rect 2183 7704 2228 7732
rect 1489 7695 1547 7701
rect 2222 7692 2228 7704
rect 2280 7692 2286 7744
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 2958 7732 2964 7744
rect 2915 7704 2964 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3881 7735 3939 7741
rect 3881 7732 3893 7735
rect 3108 7704 3893 7732
rect 3108 7692 3114 7704
rect 3881 7701 3893 7704
rect 3927 7701 3939 7735
rect 3881 7695 3939 7701
rect 1104 7642 10856 7664
rect 1104 7590 4213 7642
rect 4265 7590 4277 7642
rect 4329 7590 4341 7642
rect 4393 7590 4405 7642
rect 4457 7590 4469 7642
rect 4521 7590 7477 7642
rect 7529 7590 7541 7642
rect 7593 7590 7605 7642
rect 7657 7590 7669 7642
rect 7721 7590 7733 7642
rect 7785 7590 10856 7642
rect 1104 7568 10856 7590
rect 1857 7531 1915 7537
rect 1857 7497 1869 7531
rect 1903 7528 1915 7531
rect 1946 7528 1952 7540
rect 1903 7500 1952 7528
rect 1903 7497 1915 7500
rect 1857 7491 1915 7497
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 3050 7392 3056 7404
rect 2823 7364 3056 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 3234 7392 3240 7404
rect 3195 7364 3240 7392
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 3418 7392 3424 7404
rect 3379 7364 3424 7392
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 2593 7191 2651 7197
rect 2593 7188 2605 7191
rect 2096 7160 2605 7188
rect 2096 7148 2102 7160
rect 2593 7157 2605 7160
rect 2639 7157 2651 7191
rect 2593 7151 2651 7157
rect 3237 7191 3295 7197
rect 3237 7157 3249 7191
rect 3283 7188 3295 7191
rect 3326 7188 3332 7200
rect 3283 7160 3332 7188
rect 3283 7157 3295 7160
rect 3237 7151 3295 7157
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 1104 7098 10856 7120
rect 1104 7046 2582 7098
rect 2634 7046 2646 7098
rect 2698 7046 2710 7098
rect 2762 7046 2774 7098
rect 2826 7046 2838 7098
rect 2890 7046 5845 7098
rect 5897 7046 5909 7098
rect 5961 7046 5973 7098
rect 6025 7046 6037 7098
rect 6089 7046 6101 7098
rect 6153 7046 9109 7098
rect 9161 7046 9173 7098
rect 9225 7046 9237 7098
rect 9289 7046 9301 7098
rect 9353 7046 9365 7098
rect 9417 7046 10856 7098
rect 1104 7024 10856 7046
rect 2958 6848 2964 6860
rect 2746 6820 2964 6848
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 2746 6780 2774 6820
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 3142 6848 3148 6860
rect 3103 6820 3148 6848
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 1719 6752 2774 6780
rect 2869 6783 2927 6789
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6749 3847 6783
rect 3970 6780 3976 6792
rect 3931 6752 3976 6780
rect 3789 6743 3847 6749
rect 2884 6712 2912 6743
rect 3234 6712 3240 6724
rect 2884 6684 3240 6712
rect 3234 6672 3240 6684
rect 3292 6712 3298 6724
rect 3804 6712 3832 6743
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 3292 6684 3832 6712
rect 3292 6672 3298 6684
rect 1486 6644 1492 6656
rect 1447 6616 1492 6644
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 3878 6644 3884 6656
rect 3839 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 9950 6644 9956 6656
rect 9911 6616 9956 6644
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 1104 6554 10856 6576
rect 1104 6502 4213 6554
rect 4265 6502 4277 6554
rect 4329 6502 4341 6554
rect 4393 6502 4405 6554
rect 4457 6502 4469 6554
rect 4521 6502 7477 6554
rect 7529 6502 7541 6554
rect 7593 6502 7605 6554
rect 7657 6502 7669 6554
rect 7721 6502 7733 6554
rect 7785 6502 10856 6554
rect 1104 6480 10856 6502
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 2314 6440 2320 6452
rect 2087 6412 2320 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 2314 6400 2320 6412
rect 2372 6400 2378 6452
rect 9950 6372 9956 6384
rect 2240 6344 9956 6372
rect 2240 6313 2268 6344
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 3142 6304 3148 6316
rect 2731 6276 3148 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 2958 6236 2964 6248
rect 2919 6208 2964 6236
rect 2958 6196 2964 6208
rect 3016 6196 3022 6248
rect 4264 6236 4292 6267
rect 9950 6236 9956 6248
rect 4264 6208 9956 6236
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 1118 6128 1124 6180
rect 1176 6168 1182 6180
rect 4065 6171 4123 6177
rect 4065 6168 4077 6171
rect 1176 6140 4077 6168
rect 1176 6128 1182 6140
rect 4065 6137 4077 6140
rect 4111 6137 4123 6171
rect 4065 6131 4123 6137
rect 1104 6010 10856 6032
rect 1104 5958 2582 6010
rect 2634 5958 2646 6010
rect 2698 5958 2710 6010
rect 2762 5958 2774 6010
rect 2826 5958 2838 6010
rect 2890 5958 5845 6010
rect 5897 5958 5909 6010
rect 5961 5958 5973 6010
rect 6025 5958 6037 6010
rect 6089 5958 6101 6010
rect 6153 5958 9109 6010
rect 9161 5958 9173 6010
rect 9225 5958 9237 6010
rect 9289 5958 9301 6010
rect 9353 5958 9365 6010
rect 9417 5958 10856 6010
rect 1104 5936 10856 5958
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 4614 5896 4620 5908
rect 3283 5868 4620 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 4764 5868 4809 5896
rect 4764 5856 4770 5868
rect 1026 5720 1032 5772
rect 1084 5760 1090 5772
rect 3881 5763 3939 5769
rect 3881 5760 3893 5763
rect 1084 5732 2360 5760
rect 1084 5720 1090 5732
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 2038 5652 2044 5704
rect 2096 5692 2102 5704
rect 2332 5701 2360 5732
rect 2746 5732 3893 5760
rect 2133 5695 2191 5701
rect 2133 5692 2145 5695
rect 2096 5664 2145 5692
rect 2096 5652 2102 5664
rect 2133 5661 2145 5664
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2746 5692 2774 5732
rect 3881 5729 3893 5732
rect 3927 5729 3939 5763
rect 10965 5763 11023 5769
rect 10965 5760 10977 5763
rect 3881 5723 3939 5729
rect 4080 5732 10977 5760
rect 4080 5701 4108 5732
rect 10965 5729 10977 5732
rect 11011 5729 11023 5763
rect 10965 5723 11023 5729
rect 2363 5664 2774 5692
rect 3237 5695 3295 5701
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 3237 5661 3249 5695
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 9858 5692 9864 5704
rect 4939 5664 9864 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 3252 5624 3280 5655
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 3252 5596 9996 5624
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2130 5516 2136 5568
rect 2188 5556 2194 5568
rect 9968 5565 9996 5596
rect 2225 5559 2283 5565
rect 2225 5556 2237 5559
rect 2188 5528 2237 5556
rect 2188 5516 2194 5528
rect 2225 5525 2237 5528
rect 2271 5525 2283 5559
rect 2225 5519 2283 5525
rect 9953 5559 10011 5565
rect 9953 5525 9965 5559
rect 9999 5525 10011 5559
rect 9953 5519 10011 5525
rect 1104 5466 10856 5488
rect 1104 5414 4213 5466
rect 4265 5414 4277 5466
rect 4329 5414 4341 5466
rect 4393 5414 4405 5466
rect 4457 5414 4469 5466
rect 4521 5414 7477 5466
rect 7529 5414 7541 5466
rect 7593 5414 7605 5466
rect 7657 5414 7669 5466
rect 7721 5414 7733 5466
rect 7785 5414 10856 5466
rect 1104 5392 10856 5414
rect 3878 5352 3884 5364
rect 1688 5324 3884 5352
rect 1688 5225 1716 5324
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 9950 5352 9956 5364
rect 9911 5324 9956 5352
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 2038 5244 2044 5296
rect 2096 5284 2102 5296
rect 2590 5284 2596 5296
rect 2096 5256 2596 5284
rect 2096 5244 2102 5256
rect 2148 5225 2176 5256
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5216 2835 5219
rect 2866 5216 2872 5228
rect 2823 5188 2872 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 2332 5148 2360 5179
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5216 3019 5219
rect 3050 5216 3056 5228
rect 3007 5188 3056 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 3050 5176 3056 5188
rect 3108 5216 3114 5228
rect 3881 5219 3939 5225
rect 3881 5216 3893 5219
rect 3108 5188 3893 5216
rect 3108 5176 3114 5188
rect 3881 5185 3893 5188
rect 3927 5185 3939 5219
rect 4062 5216 4068 5228
rect 4023 5188 4068 5216
rect 3881 5179 3939 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 10134 5216 10140 5228
rect 10095 5188 10140 5216
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 4706 5148 4712 5160
rect 2332 5120 4712 5148
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 2133 5083 2191 5089
rect 2133 5049 2145 5083
rect 2179 5080 2191 5083
rect 3142 5080 3148 5092
rect 2179 5052 3148 5080
rect 2179 5049 2191 5052
rect 2133 5043 2191 5049
rect 3142 5040 3148 5052
rect 3200 5040 3206 5092
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 2777 5015 2835 5021
rect 2777 4981 2789 5015
rect 2823 5012 2835 5015
rect 2958 5012 2964 5024
rect 2823 4984 2964 5012
rect 2823 4981 2835 4984
rect 2777 4975 2835 4981
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 1104 4922 10856 4944
rect 1104 4870 2582 4922
rect 2634 4870 2646 4922
rect 2698 4870 2710 4922
rect 2762 4870 2774 4922
rect 2826 4870 2838 4922
rect 2890 4870 5845 4922
rect 5897 4870 5909 4922
rect 5961 4870 5973 4922
rect 6025 4870 6037 4922
rect 6089 4870 6101 4922
rect 6153 4870 9109 4922
rect 9161 4870 9173 4922
rect 9225 4870 9237 4922
rect 9289 4870 9301 4922
rect 9353 4870 9365 4922
rect 9417 4870 10856 4922
rect 1104 4848 10856 4870
rect 1210 4768 1216 4820
rect 1268 4808 1274 4820
rect 3050 4808 3056 4820
rect 1268 4780 3056 4808
rect 1268 4768 1274 4780
rect 3050 4768 3056 4780
rect 3108 4768 3114 4820
rect 3326 4740 3332 4752
rect 1688 4712 3332 4740
rect 1688 4613 1716 4712
rect 3326 4700 3332 4712
rect 3384 4700 3390 4752
rect 2148 4644 2544 4672
rect 2148 4613 2176 4644
rect 2516 4616 2544 4644
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 1118 4496 1124 4548
rect 1176 4536 1182 4548
rect 2332 4536 2360 4567
rect 2498 4564 2504 4616
rect 2556 4604 2562 4616
rect 2777 4607 2835 4613
rect 2777 4604 2789 4607
rect 2556 4576 2789 4604
rect 2556 4564 2562 4576
rect 2777 4573 2789 4576
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4604 3019 4607
rect 4614 4604 4620 4616
rect 3007 4576 4620 4604
rect 3007 4573 3019 4576
rect 2961 4567 3019 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 1176 4508 2360 4536
rect 1176 4496 1182 4508
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 1670 4428 1676 4480
rect 1728 4468 1734 4480
rect 2225 4471 2283 4477
rect 2225 4468 2237 4471
rect 1728 4440 2237 4468
rect 1728 4428 1734 4440
rect 2225 4437 2237 4440
rect 2271 4437 2283 4471
rect 2866 4468 2872 4480
rect 2827 4440 2872 4468
rect 2225 4431 2283 4437
rect 2866 4428 2872 4440
rect 2924 4428 2930 4480
rect 1104 4378 10856 4400
rect 1104 4326 4213 4378
rect 4265 4326 4277 4378
rect 4329 4326 4341 4378
rect 4393 4326 4405 4378
rect 4457 4326 4469 4378
rect 4521 4326 7477 4378
rect 7529 4326 7541 4378
rect 7593 4326 7605 4378
rect 7657 4326 7669 4378
rect 7721 4326 7733 4378
rect 7785 4326 10856 4378
rect 1104 4304 10856 4326
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 9953 4267 10011 4273
rect 9953 4264 9965 4267
rect 4120 4236 9965 4264
rect 4120 4224 4126 4236
rect 9953 4233 9965 4236
rect 9999 4233 10011 4267
rect 9953 4227 10011 4233
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2222 4128 2228 4140
rect 2179 4100 2228 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 1688 4060 1716 4091
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 10134 4128 10140 4140
rect 10095 4100 10140 4128
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 2866 4060 2872 4072
rect 1688 4032 2872 4060
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 2314 3924 2320 3936
rect 2275 3896 2320 3924
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 1104 3834 10856 3856
rect 1104 3782 2582 3834
rect 2634 3782 2646 3834
rect 2698 3782 2710 3834
rect 2762 3782 2774 3834
rect 2826 3782 2838 3834
rect 2890 3782 5845 3834
rect 5897 3782 5909 3834
rect 5961 3782 5973 3834
rect 6025 3782 6037 3834
rect 6089 3782 6101 3834
rect 6153 3782 9109 3834
rect 9161 3782 9173 3834
rect 9225 3782 9237 3834
rect 9289 3782 9301 3834
rect 9353 3782 9365 3834
rect 9417 3782 10856 3834
rect 1104 3760 10856 3782
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 9953 3723 10011 3729
rect 9953 3720 9965 3723
rect 9916 3692 9965 3720
rect 9916 3680 9922 3692
rect 9953 3689 9965 3692
rect 9999 3689 10011 3723
rect 9953 3683 10011 3689
rect 1670 3516 1676 3528
rect 1631 3488 1676 3516
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 1946 3476 1952 3528
rect 2004 3516 2010 3528
rect 2317 3519 2375 3525
rect 2317 3516 2329 3519
rect 2004 3488 2329 3516
rect 2004 3476 2010 3488
rect 2317 3485 2329 3488
rect 2363 3516 2375 3519
rect 9858 3516 9864 3528
rect 2363 3488 9864 3516
rect 2363 3485 2375 3488
rect 2317 3479 2375 3485
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 1489 3383 1547 3389
rect 1489 3380 1501 3383
rect 1452 3352 1501 3380
rect 1452 3340 1458 3352
rect 1489 3349 1501 3352
rect 1535 3349 1547 3383
rect 1489 3343 1547 3349
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 2133 3383 2191 3389
rect 2133 3380 2145 3383
rect 1728 3352 2145 3380
rect 1728 3340 1734 3352
rect 2133 3349 2145 3352
rect 2179 3349 2191 3383
rect 2133 3343 2191 3349
rect 1104 3290 10856 3312
rect 1104 3238 4213 3290
rect 4265 3238 4277 3290
rect 4329 3238 4341 3290
rect 4393 3238 4405 3290
rect 4457 3238 4469 3290
rect 4521 3238 7477 3290
rect 7529 3238 7541 3290
rect 7593 3238 7605 3290
rect 7657 3238 7669 3290
rect 7721 3238 7733 3290
rect 7785 3238 10856 3290
rect 1104 3216 10856 3238
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 2958 3040 2964 3052
rect 1719 3012 2964 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 9858 3040 9864 3052
rect 9819 3012 9864 3040
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 10134 2972 10140 2984
rect 10095 2944 10140 2972
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 1486 2836 1492 2848
rect 1447 2808 1492 2836
rect 1486 2796 1492 2808
rect 1544 2796 1550 2848
rect 1104 2746 10856 2768
rect 1104 2694 2582 2746
rect 2634 2694 2646 2746
rect 2698 2694 2710 2746
rect 2762 2694 2774 2746
rect 2826 2694 2838 2746
rect 2890 2694 5845 2746
rect 5897 2694 5909 2746
rect 5961 2694 5973 2746
rect 6025 2694 6037 2746
rect 6089 2694 6101 2746
rect 6153 2694 9109 2746
rect 9161 2694 9173 2746
rect 9225 2694 9237 2746
rect 9289 2694 9301 2746
rect 9353 2694 9365 2746
rect 9417 2694 10856 2746
rect 1104 2672 10856 2694
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 10965 2499 11023 2505
rect 10965 2496 10977 2499
rect 9907 2468 10977 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 10965 2465 10977 2468
rect 11011 2465 11023 2499
rect 10965 2459 11023 2465
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2130 2428 2136 2440
rect 2091 2400 2136 2428
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 2958 2428 2964 2440
rect 2915 2400 2964 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 10134 2428 10140 2440
rect 10095 2400 10140 2428
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 1394 2252 1400 2304
rect 1452 2292 1458 2304
rect 1489 2295 1547 2301
rect 1489 2292 1501 2295
rect 1452 2264 1501 2292
rect 1452 2252 1458 2264
rect 1489 2261 1501 2264
rect 1535 2261 1547 2295
rect 1489 2255 1547 2261
rect 2317 2295 2375 2301
rect 2317 2261 2329 2295
rect 2363 2292 2375 2295
rect 2774 2292 2780 2304
rect 2363 2264 2780 2292
rect 2363 2261 2375 2264
rect 2317 2255 2375 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 3050 2292 3056 2304
rect 3011 2264 3056 2292
rect 3050 2252 3056 2264
rect 3108 2252 3114 2304
rect 1104 2202 10856 2224
rect 1104 2150 4213 2202
rect 4265 2150 4277 2202
rect 4329 2150 4341 2202
rect 4393 2150 4405 2202
rect 4457 2150 4469 2202
rect 4521 2150 7477 2202
rect 7529 2150 7541 2202
rect 7593 2150 7605 2202
rect 7657 2150 7669 2202
rect 7721 2150 7733 2202
rect 7785 2150 10856 2202
rect 1104 2128 10856 2150
<< via1 >>
rect 10968 78659 11020 78668
rect 10968 78625 10977 78659
rect 10977 78625 11011 78659
rect 11011 78625 11020 78659
rect 10968 78616 11020 78625
rect 2582 77766 2634 77818
rect 2646 77766 2698 77818
rect 2710 77766 2762 77818
rect 2774 77766 2826 77818
rect 2838 77766 2890 77818
rect 5845 77766 5897 77818
rect 5909 77766 5961 77818
rect 5973 77766 6025 77818
rect 6037 77766 6089 77818
rect 6101 77766 6153 77818
rect 9109 77766 9161 77818
rect 9173 77766 9225 77818
rect 9237 77766 9289 77818
rect 9301 77766 9353 77818
rect 9365 77766 9417 77818
rect 9496 77664 9548 77716
rect 1768 77596 1820 77648
rect 1400 77503 1452 77512
rect 1400 77469 1409 77503
rect 1409 77469 1443 77503
rect 1443 77469 1452 77503
rect 1400 77460 1452 77469
rect 2044 77503 2096 77512
rect 2044 77469 2053 77503
rect 2053 77469 2087 77503
rect 2087 77469 2096 77503
rect 2044 77460 2096 77469
rect 2964 77460 3016 77512
rect 3792 77503 3844 77512
rect 3792 77469 3801 77503
rect 3801 77469 3835 77503
rect 3835 77469 3844 77503
rect 3792 77460 3844 77469
rect 5540 77460 5592 77512
rect 1676 77324 1728 77376
rect 2504 77324 2556 77376
rect 3976 77367 4028 77376
rect 3976 77333 3985 77367
rect 3985 77333 4019 77367
rect 4019 77333 4028 77367
rect 3976 77324 4028 77333
rect 10048 77367 10100 77376
rect 10048 77333 10057 77367
rect 10057 77333 10091 77367
rect 10091 77333 10100 77367
rect 10048 77324 10100 77333
rect 4213 77222 4265 77274
rect 4277 77222 4329 77274
rect 4341 77222 4393 77274
rect 4405 77222 4457 77274
rect 4469 77222 4521 77274
rect 7477 77222 7529 77274
rect 7541 77222 7593 77274
rect 7605 77222 7657 77274
rect 7669 77222 7721 77274
rect 7733 77222 7785 77274
rect 9588 77120 9640 77172
rect 1308 76984 1360 77036
rect 1492 76984 1544 77036
rect 3056 76984 3108 77036
rect 8300 76984 8352 77036
rect 9680 76984 9732 77036
rect 1584 76823 1636 76832
rect 1584 76789 1593 76823
rect 1593 76789 1627 76823
rect 1627 76789 1636 76823
rect 1584 76780 1636 76789
rect 2228 76823 2280 76832
rect 2228 76789 2237 76823
rect 2237 76789 2271 76823
rect 2271 76789 2280 76823
rect 2228 76780 2280 76789
rect 3608 76780 3660 76832
rect 10048 76823 10100 76832
rect 10048 76789 10057 76823
rect 10057 76789 10091 76823
rect 10091 76789 10100 76823
rect 10048 76780 10100 76789
rect 2582 76678 2634 76730
rect 2646 76678 2698 76730
rect 2710 76678 2762 76730
rect 2774 76678 2826 76730
rect 2838 76678 2890 76730
rect 5845 76678 5897 76730
rect 5909 76678 5961 76730
rect 5973 76678 6025 76730
rect 6037 76678 6089 76730
rect 6101 76678 6153 76730
rect 9109 76678 9161 76730
rect 9173 76678 9225 76730
rect 9237 76678 9289 76730
rect 9301 76678 9353 76730
rect 9365 76678 9417 76730
rect 1400 76415 1452 76424
rect 1400 76381 1409 76415
rect 1409 76381 1443 76415
rect 1443 76381 1452 76415
rect 1400 76372 1452 76381
rect 9772 76372 9824 76424
rect 1492 76236 1544 76288
rect 4213 76134 4265 76186
rect 4277 76134 4329 76186
rect 4341 76134 4393 76186
rect 4405 76134 4457 76186
rect 4469 76134 4521 76186
rect 7477 76134 7529 76186
rect 7541 76134 7593 76186
rect 7605 76134 7657 76186
rect 7669 76134 7721 76186
rect 7733 76134 7785 76186
rect 3056 76032 3108 76084
rect 1308 75896 1360 75948
rect 6276 75828 6328 75880
rect 10048 75735 10100 75744
rect 10048 75701 10057 75735
rect 10057 75701 10091 75735
rect 10091 75701 10100 75735
rect 10048 75692 10100 75701
rect 2582 75590 2634 75642
rect 2646 75590 2698 75642
rect 2710 75590 2762 75642
rect 2774 75590 2826 75642
rect 2838 75590 2890 75642
rect 5845 75590 5897 75642
rect 5909 75590 5961 75642
rect 5973 75590 6025 75642
rect 6037 75590 6089 75642
rect 6101 75590 6153 75642
rect 9109 75590 9161 75642
rect 9173 75590 9225 75642
rect 9237 75590 9289 75642
rect 9301 75590 9353 75642
rect 9365 75590 9417 75642
rect 3148 75420 3200 75472
rect 1400 75327 1452 75336
rect 1400 75293 1409 75327
rect 1409 75293 1443 75327
rect 1443 75293 1452 75327
rect 1400 75284 1452 75293
rect 2044 75327 2096 75336
rect 2044 75293 2053 75327
rect 2053 75293 2087 75327
rect 2087 75293 2096 75327
rect 2044 75284 2096 75293
rect 9864 75327 9916 75336
rect 9864 75293 9873 75327
rect 9873 75293 9907 75327
rect 9907 75293 9916 75327
rect 9864 75284 9916 75293
rect 2964 75148 3016 75200
rect 10048 75191 10100 75200
rect 10048 75157 10057 75191
rect 10057 75157 10091 75191
rect 10091 75157 10100 75191
rect 10048 75148 10100 75157
rect 4213 75046 4265 75098
rect 4277 75046 4329 75098
rect 4341 75046 4393 75098
rect 4405 75046 4457 75098
rect 4469 75046 4521 75098
rect 7477 75046 7529 75098
rect 7541 75046 7593 75098
rect 7605 75046 7657 75098
rect 7669 75046 7721 75098
rect 7733 75046 7785 75098
rect 1676 74919 1728 74928
rect 1676 74885 1685 74919
rect 1685 74885 1719 74919
rect 1719 74885 1728 74919
rect 1676 74876 1728 74885
rect 2228 74876 2280 74928
rect 5540 74944 5592 74996
rect 6552 74876 6604 74928
rect 2136 74808 2188 74860
rect 2596 74851 2648 74860
rect 1676 74740 1728 74792
rect 2596 74817 2605 74851
rect 2605 74817 2639 74851
rect 2639 74817 2648 74851
rect 2596 74808 2648 74817
rect 3700 74808 3752 74860
rect 3516 74740 3568 74792
rect 1124 74672 1176 74724
rect 2596 74672 2648 74724
rect 6276 74604 6328 74656
rect 2582 74502 2634 74554
rect 2646 74502 2698 74554
rect 2710 74502 2762 74554
rect 2774 74502 2826 74554
rect 2838 74502 2890 74554
rect 5845 74502 5897 74554
rect 5909 74502 5961 74554
rect 5973 74502 6025 74554
rect 6037 74502 6089 74554
rect 6101 74502 6153 74554
rect 9109 74502 9161 74554
rect 9173 74502 9225 74554
rect 9237 74502 9289 74554
rect 9301 74502 9353 74554
rect 9365 74502 9417 74554
rect 9864 74400 9916 74452
rect 9680 74332 9732 74384
rect 1584 74264 1636 74316
rect 2136 74196 2188 74248
rect 2688 74239 2740 74248
rect 1584 74171 1636 74180
rect 1584 74137 1593 74171
rect 1593 74137 1627 74171
rect 1627 74137 1636 74171
rect 1584 74128 1636 74137
rect 2688 74205 2697 74239
rect 2697 74205 2731 74239
rect 2731 74205 2740 74239
rect 2688 74196 2740 74205
rect 2780 74239 2832 74248
rect 2780 74205 2789 74239
rect 2789 74205 2823 74239
rect 2823 74205 2832 74239
rect 2780 74196 2832 74205
rect 3332 74128 3384 74180
rect 1676 74060 1728 74112
rect 2504 74060 2556 74112
rect 5632 74264 5684 74316
rect 3792 74239 3844 74248
rect 3792 74205 3801 74239
rect 3801 74205 3835 74239
rect 3835 74205 3844 74239
rect 3792 74196 3844 74205
rect 3976 74196 4028 74248
rect 4804 74196 4856 74248
rect 9864 74239 9916 74248
rect 9864 74205 9873 74239
rect 9873 74205 9907 74239
rect 9907 74205 9916 74239
rect 9864 74196 9916 74205
rect 3700 74128 3752 74180
rect 4988 74128 5040 74180
rect 4068 74060 4120 74112
rect 10048 74103 10100 74112
rect 10048 74069 10057 74103
rect 10057 74069 10091 74103
rect 10091 74069 10100 74103
rect 10048 74060 10100 74069
rect 4213 73958 4265 74010
rect 4277 73958 4329 74010
rect 4341 73958 4393 74010
rect 4405 73958 4457 74010
rect 4469 73958 4521 74010
rect 7477 73958 7529 74010
rect 7541 73958 7593 74010
rect 7605 73958 7657 74010
rect 7669 73958 7721 74010
rect 7733 73958 7785 74010
rect 2504 73856 2556 73908
rect 1492 73788 1544 73840
rect 2964 73788 3016 73840
rect 3608 73788 3660 73840
rect 2136 73720 2188 73772
rect 2412 73720 2464 73772
rect 3516 73763 3568 73772
rect 3516 73729 3525 73763
rect 3525 73729 3559 73763
rect 3559 73729 3568 73763
rect 3516 73720 3568 73729
rect 1492 73584 1544 73636
rect 1676 73584 1728 73636
rect 480 73516 532 73568
rect 2780 73652 2832 73704
rect 2964 73652 3016 73704
rect 3792 73652 3844 73704
rect 4712 73831 4764 73840
rect 4712 73797 4721 73831
rect 4721 73797 4755 73831
rect 4755 73797 4764 73831
rect 8300 73856 8352 73908
rect 4712 73788 4764 73797
rect 9772 73788 9824 73840
rect 4528 73763 4580 73772
rect 4528 73729 4557 73763
rect 4557 73729 4580 73763
rect 4528 73720 4580 73729
rect 4804 73763 4856 73772
rect 4804 73729 4809 73763
rect 4809 73729 4843 73763
rect 4843 73729 4856 73763
rect 4804 73720 4856 73729
rect 4988 73720 5040 73772
rect 4988 73584 5040 73636
rect 9864 73516 9916 73568
rect 10048 73559 10100 73568
rect 10048 73525 10057 73559
rect 10057 73525 10091 73559
rect 10091 73525 10100 73559
rect 10048 73516 10100 73525
rect 2582 73414 2634 73466
rect 2646 73414 2698 73466
rect 2710 73414 2762 73466
rect 2774 73414 2826 73466
rect 2838 73414 2890 73466
rect 5845 73414 5897 73466
rect 5909 73414 5961 73466
rect 5973 73414 6025 73466
rect 6037 73414 6089 73466
rect 6101 73414 6153 73466
rect 9109 73414 9161 73466
rect 9173 73414 9225 73466
rect 9237 73414 9289 73466
rect 9301 73414 9353 73466
rect 9365 73414 9417 73466
rect 1584 73312 1636 73364
rect 4804 73312 4856 73364
rect 1492 73108 1544 73160
rect 1676 73151 1728 73160
rect 1676 73117 1685 73151
rect 1685 73117 1719 73151
rect 1719 73117 1728 73151
rect 1676 73108 1728 73117
rect 2136 73108 2188 73160
rect 2412 73108 2464 73160
rect 2872 73151 2924 73160
rect 2872 73117 2881 73151
rect 2881 73117 2915 73151
rect 2915 73117 2924 73151
rect 2872 73108 2924 73117
rect 2964 73108 3016 73160
rect 3516 73176 3568 73228
rect 4528 73176 4580 73228
rect 1584 73083 1636 73092
rect 1584 73049 1593 73083
rect 1593 73049 1627 73083
rect 1627 73049 1636 73083
rect 1584 73040 1636 73049
rect 848 72972 900 73024
rect 10048 73015 10100 73024
rect 10048 72981 10057 73015
rect 10057 72981 10091 73015
rect 10091 72981 10100 73015
rect 10048 72972 10100 72981
rect 4213 72870 4265 72922
rect 4277 72870 4329 72922
rect 4341 72870 4393 72922
rect 4405 72870 4457 72922
rect 4469 72870 4521 72922
rect 7477 72870 7529 72922
rect 7541 72870 7593 72922
rect 7605 72870 7657 72922
rect 7669 72870 7721 72922
rect 7733 72870 7785 72922
rect 1492 72700 1544 72752
rect 1400 72675 1452 72684
rect 1400 72641 1409 72675
rect 1409 72641 1443 72675
rect 1443 72641 1452 72675
rect 1400 72632 1452 72641
rect 2044 72675 2096 72684
rect 2044 72641 2053 72675
rect 2053 72641 2087 72675
rect 2087 72641 2096 72675
rect 2044 72632 2096 72641
rect 2136 72632 2188 72684
rect 1584 72564 1636 72616
rect 3792 72564 3844 72616
rect 3976 72607 4028 72616
rect 3976 72573 3985 72607
rect 3985 72573 4019 72607
rect 4019 72573 4028 72607
rect 3976 72564 4028 72573
rect 7012 72496 7064 72548
rect 1676 72428 1728 72480
rect 2320 72428 2372 72480
rect 2504 72428 2556 72480
rect 5724 72428 5776 72480
rect 2582 72326 2634 72378
rect 2646 72326 2698 72378
rect 2710 72326 2762 72378
rect 2774 72326 2826 72378
rect 2838 72326 2890 72378
rect 5845 72326 5897 72378
rect 5909 72326 5961 72378
rect 5973 72326 6025 72378
rect 6037 72326 6089 72378
rect 6101 72326 6153 72378
rect 9109 72326 9161 72378
rect 9173 72326 9225 72378
rect 9237 72326 9289 72378
rect 9301 72326 9353 72378
rect 9365 72326 9417 72378
rect 3608 72224 3660 72276
rect 2504 72156 2556 72208
rect 1400 72063 1452 72072
rect 1400 72029 1409 72063
rect 1409 72029 1443 72063
rect 1443 72029 1452 72063
rect 1400 72020 1452 72029
rect 2412 72020 2464 72072
rect 3148 72088 3200 72140
rect 2964 72020 3016 72072
rect 3884 72020 3936 72072
rect 4068 72063 4120 72072
rect 4068 72029 4077 72063
rect 4077 72029 4111 72063
rect 4111 72029 4120 72063
rect 4068 72020 4120 72029
rect 6460 71952 6512 72004
rect 2872 71884 2924 71936
rect 9864 71884 9916 71936
rect 10048 71927 10100 71936
rect 10048 71893 10057 71927
rect 10057 71893 10091 71927
rect 10091 71893 10100 71927
rect 10048 71884 10100 71893
rect 4213 71782 4265 71834
rect 4277 71782 4329 71834
rect 4341 71782 4393 71834
rect 4405 71782 4457 71834
rect 4469 71782 4521 71834
rect 7477 71782 7529 71834
rect 7541 71782 7593 71834
rect 7605 71782 7657 71834
rect 7669 71782 7721 71834
rect 7733 71782 7785 71834
rect 1400 71587 1452 71596
rect 1400 71553 1409 71587
rect 1409 71553 1443 71587
rect 1443 71553 1452 71587
rect 1400 71544 1452 71553
rect 4620 71680 4672 71732
rect 2320 71655 2372 71664
rect 2320 71621 2329 71655
rect 2329 71621 2363 71655
rect 2363 71621 2372 71655
rect 2320 71612 2372 71621
rect 2964 71544 3016 71596
rect 3792 71544 3844 71596
rect 9864 71587 9916 71596
rect 9864 71553 9873 71587
rect 9873 71553 9907 71587
rect 9907 71553 9916 71587
rect 9864 71544 9916 71553
rect 2872 71476 2924 71528
rect 2504 71340 2556 71392
rect 9864 71340 9916 71392
rect 10048 71383 10100 71392
rect 10048 71349 10057 71383
rect 10057 71349 10091 71383
rect 10091 71349 10100 71383
rect 10048 71340 10100 71349
rect 2582 71238 2634 71290
rect 2646 71238 2698 71290
rect 2710 71238 2762 71290
rect 2774 71238 2826 71290
rect 2838 71238 2890 71290
rect 5845 71238 5897 71290
rect 5909 71238 5961 71290
rect 5973 71238 6025 71290
rect 6037 71238 6089 71290
rect 6101 71238 6153 71290
rect 9109 71238 9161 71290
rect 9173 71238 9225 71290
rect 9237 71238 9289 71290
rect 9301 71238 9353 71290
rect 9365 71238 9417 71290
rect 3976 71000 4028 71052
rect 1400 70975 1452 70984
rect 1400 70941 1409 70975
rect 1409 70941 1443 70975
rect 1443 70941 1452 70975
rect 1400 70932 1452 70941
rect 3884 70932 3936 70984
rect 2412 70796 2464 70848
rect 3700 70796 3752 70848
rect 3884 70796 3936 70848
rect 4213 70694 4265 70746
rect 4277 70694 4329 70746
rect 4341 70694 4393 70746
rect 4405 70694 4457 70746
rect 4469 70694 4521 70746
rect 7477 70694 7529 70746
rect 7541 70694 7593 70746
rect 7605 70694 7657 70746
rect 7669 70694 7721 70746
rect 7733 70694 7785 70746
rect 2044 70592 2096 70644
rect 10692 70592 10744 70644
rect 1400 70499 1452 70508
rect 1400 70465 1409 70499
rect 1409 70465 1443 70499
rect 1443 70465 1452 70499
rect 1400 70456 1452 70465
rect 9864 70499 9916 70508
rect 9864 70465 9873 70499
rect 9873 70465 9907 70499
rect 9907 70465 9916 70499
rect 9864 70456 9916 70465
rect 2582 70150 2634 70202
rect 2646 70150 2698 70202
rect 2710 70150 2762 70202
rect 2774 70150 2826 70202
rect 2838 70150 2890 70202
rect 5845 70150 5897 70202
rect 5909 70150 5961 70202
rect 5973 70150 6025 70202
rect 6037 70150 6089 70202
rect 6101 70150 6153 70202
rect 9109 70150 9161 70202
rect 9173 70150 9225 70202
rect 9237 70150 9289 70202
rect 9301 70150 9353 70202
rect 9365 70150 9417 70202
rect 1400 69887 1452 69896
rect 1400 69853 1409 69887
rect 1409 69853 1443 69887
rect 1443 69853 1452 69887
rect 1400 69844 1452 69853
rect 2320 69708 2372 69760
rect 10048 69751 10100 69760
rect 10048 69717 10057 69751
rect 10057 69717 10091 69751
rect 10091 69717 10100 69751
rect 10048 69708 10100 69717
rect 4213 69606 4265 69658
rect 4277 69606 4329 69658
rect 4341 69606 4393 69658
rect 4405 69606 4457 69658
rect 4469 69606 4521 69658
rect 7477 69606 7529 69658
rect 7541 69606 7593 69658
rect 7605 69606 7657 69658
rect 7669 69606 7721 69658
rect 7733 69606 7785 69658
rect 1400 69411 1452 69420
rect 1400 69377 1409 69411
rect 1409 69377 1443 69411
rect 1443 69377 1452 69411
rect 1400 69368 1452 69377
rect 1768 69164 1820 69216
rect 10048 69207 10100 69216
rect 10048 69173 10057 69207
rect 10057 69173 10091 69207
rect 10091 69173 10100 69207
rect 10048 69164 10100 69173
rect 2582 69062 2634 69114
rect 2646 69062 2698 69114
rect 2710 69062 2762 69114
rect 2774 69062 2826 69114
rect 2838 69062 2890 69114
rect 5845 69062 5897 69114
rect 5909 69062 5961 69114
rect 5973 69062 6025 69114
rect 6037 69062 6089 69114
rect 6101 69062 6153 69114
rect 9109 69062 9161 69114
rect 9173 69062 9225 69114
rect 9237 69062 9289 69114
rect 9301 69062 9353 69114
rect 9365 69062 9417 69114
rect 3332 68960 3384 69012
rect 6184 68960 6236 69012
rect 1400 68799 1452 68808
rect 1400 68765 1409 68799
rect 1409 68765 1443 68799
rect 1443 68765 1452 68799
rect 1400 68756 1452 68765
rect 1492 68620 1544 68672
rect 4213 68518 4265 68570
rect 4277 68518 4329 68570
rect 4341 68518 4393 68570
rect 4405 68518 4457 68570
rect 4469 68518 4521 68570
rect 7477 68518 7529 68570
rect 7541 68518 7593 68570
rect 7605 68518 7657 68570
rect 7669 68518 7721 68570
rect 7733 68518 7785 68570
rect 1400 68323 1452 68332
rect 1400 68289 1409 68323
rect 1409 68289 1443 68323
rect 1443 68289 1452 68323
rect 1400 68280 1452 68289
rect 9864 68323 9916 68332
rect 9864 68289 9873 68323
rect 9873 68289 9907 68323
rect 9907 68289 9916 68323
rect 9864 68280 9916 68289
rect 10048 68187 10100 68196
rect 10048 68153 10057 68187
rect 10057 68153 10091 68187
rect 10091 68153 10100 68187
rect 10048 68144 10100 68153
rect 1860 68076 1912 68128
rect 2582 67974 2634 68026
rect 2646 67974 2698 68026
rect 2710 67974 2762 68026
rect 2774 67974 2826 68026
rect 2838 67974 2890 68026
rect 5845 67974 5897 68026
rect 5909 67974 5961 68026
rect 5973 67974 6025 68026
rect 6037 67974 6089 68026
rect 6101 67974 6153 68026
rect 9109 67974 9161 68026
rect 9173 67974 9225 68026
rect 9237 67974 9289 68026
rect 9301 67974 9353 68026
rect 9365 67974 9417 68026
rect 2136 67872 2188 67924
rect 1952 67804 2004 67856
rect 1400 67711 1452 67720
rect 1400 67677 1409 67711
rect 1409 67677 1443 67711
rect 1443 67677 1452 67711
rect 1400 67668 1452 67677
rect 2228 67711 2280 67720
rect 2228 67677 2237 67711
rect 2237 67677 2271 67711
rect 2271 67677 2280 67711
rect 2228 67668 2280 67677
rect 9772 67668 9824 67720
rect 10048 67575 10100 67584
rect 10048 67541 10057 67575
rect 10057 67541 10091 67575
rect 10091 67541 10100 67575
rect 10048 67532 10100 67541
rect 4213 67430 4265 67482
rect 4277 67430 4329 67482
rect 4341 67430 4393 67482
rect 4405 67430 4457 67482
rect 4469 67430 4521 67482
rect 7477 67430 7529 67482
rect 7541 67430 7593 67482
rect 7605 67430 7657 67482
rect 7669 67430 7721 67482
rect 7733 67430 7785 67482
rect 1216 67192 1268 67244
rect 2228 67235 2280 67244
rect 2228 67201 2237 67235
rect 2237 67201 2271 67235
rect 2271 67201 2280 67235
rect 2228 67192 2280 67201
rect 9588 67192 9640 67244
rect 2320 67124 2372 67176
rect 3056 67124 3108 67176
rect 1584 67031 1636 67040
rect 1584 66997 1593 67031
rect 1593 66997 1627 67031
rect 1627 66997 1636 67031
rect 1584 66988 1636 66997
rect 2320 66988 2372 67040
rect 3516 66988 3568 67040
rect 4068 66988 4120 67040
rect 10048 67031 10100 67040
rect 10048 66997 10057 67031
rect 10057 66997 10091 67031
rect 10091 66997 10100 67031
rect 10048 66988 10100 66997
rect 2582 66886 2634 66938
rect 2646 66886 2698 66938
rect 2710 66886 2762 66938
rect 2774 66886 2826 66938
rect 2838 66886 2890 66938
rect 5845 66886 5897 66938
rect 5909 66886 5961 66938
rect 5973 66886 6025 66938
rect 6037 66886 6089 66938
rect 6101 66886 6153 66938
rect 9109 66886 9161 66938
rect 9173 66886 9225 66938
rect 9237 66886 9289 66938
rect 9301 66886 9353 66938
rect 9365 66886 9417 66938
rect 9864 66784 9916 66836
rect 2412 66716 2464 66768
rect 2688 66716 2740 66768
rect 1308 66580 1360 66632
rect 2228 66580 2280 66632
rect 2504 66580 2556 66632
rect 2872 66580 2924 66632
rect 3516 66580 3568 66632
rect 3792 66580 3844 66632
rect 2412 66444 2464 66496
rect 4213 66342 4265 66394
rect 4277 66342 4329 66394
rect 4341 66342 4393 66394
rect 4405 66342 4457 66394
rect 4469 66342 4521 66394
rect 7477 66342 7529 66394
rect 7541 66342 7593 66394
rect 7605 66342 7657 66394
rect 7669 66342 7721 66394
rect 7733 66342 7785 66394
rect 2228 66240 2280 66292
rect 1676 66215 1728 66224
rect 1676 66181 1685 66215
rect 1685 66181 1719 66215
rect 1719 66181 1728 66215
rect 1676 66172 1728 66181
rect 2872 66240 2924 66292
rect 3700 66215 3752 66224
rect 756 66036 808 66088
rect 2504 66104 2556 66156
rect 2688 66147 2740 66156
rect 2688 66113 2697 66147
rect 2697 66113 2731 66147
rect 2731 66113 2740 66147
rect 2688 66104 2740 66113
rect 2872 66104 2924 66156
rect 3700 66181 3709 66215
rect 3709 66181 3743 66215
rect 3743 66181 3752 66215
rect 3700 66172 3752 66181
rect 3608 66147 3660 66156
rect 3608 66113 3617 66147
rect 3617 66113 3651 66147
rect 3651 66113 3660 66147
rect 3608 66104 3660 66113
rect 3976 66104 4028 66156
rect 9680 66104 9732 66156
rect 9772 66036 9824 66088
rect 10048 65943 10100 65952
rect 10048 65909 10057 65943
rect 10057 65909 10091 65943
rect 10091 65909 10100 65943
rect 10048 65900 10100 65909
rect 2582 65798 2634 65850
rect 2646 65798 2698 65850
rect 2710 65798 2762 65850
rect 2774 65798 2826 65850
rect 2838 65798 2890 65850
rect 5845 65798 5897 65850
rect 5909 65798 5961 65850
rect 5973 65798 6025 65850
rect 6037 65798 6089 65850
rect 6101 65798 6153 65850
rect 9109 65798 9161 65850
rect 9173 65798 9225 65850
rect 9237 65798 9289 65850
rect 9301 65798 9353 65850
rect 9365 65798 9417 65850
rect 1032 65356 1084 65408
rect 3608 65696 3660 65748
rect 3792 65628 3844 65680
rect 2228 65560 2280 65612
rect 3240 65603 3292 65612
rect 3240 65569 3249 65603
rect 3249 65569 3283 65603
rect 3283 65569 3292 65603
rect 3240 65560 3292 65569
rect 3976 65560 4028 65612
rect 1400 65535 1452 65544
rect 1400 65501 1409 65535
rect 1409 65501 1443 65535
rect 1443 65501 1452 65535
rect 1400 65492 1452 65501
rect 3516 65492 3568 65544
rect 9864 65535 9916 65544
rect 9864 65501 9873 65535
rect 9873 65501 9907 65535
rect 9907 65501 9916 65535
rect 9864 65492 9916 65501
rect 1676 65356 1728 65408
rect 10048 65399 10100 65408
rect 10048 65365 10057 65399
rect 10057 65365 10091 65399
rect 10091 65365 10100 65399
rect 10048 65356 10100 65365
rect 4213 65254 4265 65306
rect 4277 65254 4329 65306
rect 4341 65254 4393 65306
rect 4405 65254 4457 65306
rect 4469 65254 4521 65306
rect 7477 65254 7529 65306
rect 7541 65254 7593 65306
rect 7605 65254 7657 65306
rect 7669 65254 7721 65306
rect 7733 65254 7785 65306
rect 848 65152 900 65204
rect 1216 65152 1268 65204
rect 9588 65152 9640 65204
rect 2044 65084 2096 65136
rect 1308 65016 1360 65068
rect 2228 65016 2280 65068
rect 5356 65084 5408 65136
rect 2964 65016 3016 65068
rect 2504 64948 2556 65000
rect 6644 64948 6696 65000
rect 2228 64880 2280 64932
rect 2582 64710 2634 64762
rect 2646 64710 2698 64762
rect 2710 64710 2762 64762
rect 2774 64710 2826 64762
rect 2838 64710 2890 64762
rect 5845 64710 5897 64762
rect 5909 64710 5961 64762
rect 5973 64710 6025 64762
rect 6037 64710 6089 64762
rect 6101 64710 6153 64762
rect 9109 64710 9161 64762
rect 9173 64710 9225 64762
rect 9237 64710 9289 64762
rect 9301 64710 9353 64762
rect 9365 64710 9417 64762
rect 9864 64540 9916 64592
rect 1400 64404 1452 64456
rect 1768 64447 1820 64456
rect 1768 64413 1777 64447
rect 1777 64413 1811 64447
rect 1811 64413 1820 64447
rect 1768 64404 1820 64413
rect 2964 64472 3016 64524
rect 2780 64404 2832 64456
rect 2872 64404 2924 64456
rect 3056 64404 3108 64456
rect 9772 64404 9824 64456
rect 7196 64336 7248 64388
rect 10048 64311 10100 64320
rect 10048 64277 10057 64311
rect 10057 64277 10091 64311
rect 10091 64277 10100 64311
rect 10048 64268 10100 64277
rect 4213 64166 4265 64218
rect 4277 64166 4329 64218
rect 4341 64166 4393 64218
rect 4405 64166 4457 64218
rect 4469 64166 4521 64218
rect 7477 64166 7529 64218
rect 7541 64166 7593 64218
rect 7605 64166 7657 64218
rect 7669 64166 7721 64218
rect 7733 64166 7785 64218
rect 1492 64064 1544 64116
rect 9680 64064 9732 64116
rect 8392 63996 8444 64048
rect 1492 63971 1544 63980
rect 1492 63937 1501 63971
rect 1501 63937 1535 63971
rect 1535 63937 1544 63971
rect 1492 63928 1544 63937
rect 2504 63971 2556 63980
rect 2504 63937 2513 63971
rect 2513 63937 2547 63971
rect 2547 63937 2556 63971
rect 2504 63928 2556 63937
rect 2780 63971 2832 63980
rect 2780 63937 2789 63971
rect 2789 63937 2823 63971
rect 2823 63937 2832 63971
rect 2780 63928 2832 63937
rect 2964 63928 3016 63980
rect 9864 63971 9916 63980
rect 9864 63937 9873 63971
rect 9873 63937 9907 63971
rect 9907 63937 9916 63971
rect 9864 63928 9916 63937
rect 9772 63792 9824 63844
rect 8300 63724 8352 63776
rect 10048 63767 10100 63776
rect 10048 63733 10057 63767
rect 10057 63733 10091 63767
rect 10091 63733 10100 63767
rect 10048 63724 10100 63733
rect 2582 63622 2634 63674
rect 2646 63622 2698 63674
rect 2710 63622 2762 63674
rect 2774 63622 2826 63674
rect 2838 63622 2890 63674
rect 5845 63622 5897 63674
rect 5909 63622 5961 63674
rect 5973 63622 6025 63674
rect 6037 63622 6089 63674
rect 6101 63622 6153 63674
rect 9109 63622 9161 63674
rect 9173 63622 9225 63674
rect 9237 63622 9289 63674
rect 9301 63622 9353 63674
rect 9365 63622 9417 63674
rect 1768 63520 1820 63572
rect 2044 63520 2096 63572
rect 2320 63520 2372 63572
rect 2504 63520 2556 63572
rect 9864 63452 9916 63504
rect 2872 63384 2924 63436
rect 3332 63384 3384 63436
rect 3516 63384 3568 63436
rect 1492 63316 1544 63368
rect 1860 63359 1912 63368
rect 1860 63325 1869 63359
rect 1869 63325 1903 63359
rect 1903 63325 1912 63359
rect 1860 63316 1912 63325
rect 2044 63316 2096 63368
rect 2780 63359 2832 63368
rect 2780 63325 2789 63359
rect 2789 63325 2823 63359
rect 2823 63325 2832 63359
rect 3976 63359 4028 63368
rect 2780 63316 2832 63325
rect 3976 63325 3985 63359
rect 3985 63325 4019 63359
rect 4019 63325 4028 63359
rect 3976 63316 4028 63325
rect 9864 63359 9916 63368
rect 9864 63325 9873 63359
rect 9873 63325 9907 63359
rect 9907 63325 9916 63359
rect 9864 63316 9916 63325
rect 6920 63248 6972 63300
rect 2596 63223 2648 63232
rect 2596 63189 2605 63223
rect 2605 63189 2639 63223
rect 2639 63189 2648 63223
rect 2596 63180 2648 63189
rect 2688 63180 2740 63232
rect 10048 63223 10100 63232
rect 10048 63189 10057 63223
rect 10057 63189 10091 63223
rect 10091 63189 10100 63223
rect 10048 63180 10100 63189
rect 4213 63078 4265 63130
rect 4277 63078 4329 63130
rect 4341 63078 4393 63130
rect 4405 63078 4457 63130
rect 4469 63078 4521 63130
rect 7477 63078 7529 63130
rect 7541 63078 7593 63130
rect 7605 63078 7657 63130
rect 7669 63078 7721 63130
rect 7733 63078 7785 63130
rect 2964 62976 3016 63028
rect 1492 62840 1544 62892
rect 1768 62840 1820 62892
rect 1952 62883 2004 62892
rect 1952 62849 1961 62883
rect 1961 62849 1995 62883
rect 1995 62849 2004 62883
rect 1952 62840 2004 62849
rect 2044 62883 2096 62892
rect 2044 62849 2053 62883
rect 2053 62849 2087 62883
rect 2087 62849 2096 62883
rect 2044 62840 2096 62849
rect 2872 62840 2924 62892
rect 2596 62772 2648 62824
rect 1952 62704 2004 62756
rect 2044 62704 2096 62756
rect 2688 62704 2740 62756
rect 8484 62704 8536 62756
rect 9864 62636 9916 62688
rect 2582 62534 2634 62586
rect 2646 62534 2698 62586
rect 2710 62534 2762 62586
rect 2774 62534 2826 62586
rect 2838 62534 2890 62586
rect 5845 62534 5897 62586
rect 5909 62534 5961 62586
rect 5973 62534 6025 62586
rect 6037 62534 6089 62586
rect 6101 62534 6153 62586
rect 9109 62534 9161 62586
rect 9173 62534 9225 62586
rect 9237 62534 9289 62586
rect 9301 62534 9353 62586
rect 9365 62534 9417 62586
rect 2044 62432 2096 62484
rect 2412 62432 2464 62484
rect 1768 62296 1820 62348
rect 3240 62339 3292 62348
rect 3240 62305 3249 62339
rect 3249 62305 3283 62339
rect 3283 62305 3292 62339
rect 3240 62296 3292 62305
rect 3792 62160 3844 62212
rect 1492 62135 1544 62144
rect 1492 62101 1501 62135
rect 1501 62101 1535 62135
rect 1535 62101 1544 62135
rect 1492 62092 1544 62101
rect 1952 62092 2004 62144
rect 2136 62092 2188 62144
rect 10048 62135 10100 62144
rect 10048 62101 10057 62135
rect 10057 62101 10091 62135
rect 10091 62101 10100 62135
rect 10048 62092 10100 62101
rect 4213 61990 4265 62042
rect 4277 61990 4329 62042
rect 4341 61990 4393 62042
rect 4405 61990 4457 62042
rect 4469 61990 4521 62042
rect 7477 61990 7529 62042
rect 7541 61990 7593 62042
rect 7605 61990 7657 62042
rect 7669 61990 7721 62042
rect 7733 61990 7785 62042
rect 2320 61795 2372 61804
rect 2320 61761 2329 61795
rect 2329 61761 2363 61795
rect 2363 61761 2372 61795
rect 2320 61752 2372 61761
rect 3700 61684 3752 61736
rect 1400 61548 1452 61600
rect 1768 61548 1820 61600
rect 10048 61591 10100 61600
rect 10048 61557 10057 61591
rect 10057 61557 10091 61591
rect 10091 61557 10100 61591
rect 10048 61548 10100 61557
rect 2582 61446 2634 61498
rect 2646 61446 2698 61498
rect 2710 61446 2762 61498
rect 2774 61446 2826 61498
rect 2838 61446 2890 61498
rect 5845 61446 5897 61498
rect 5909 61446 5961 61498
rect 5973 61446 6025 61498
rect 6037 61446 6089 61498
rect 6101 61446 6153 61498
rect 9109 61446 9161 61498
rect 9173 61446 9225 61498
rect 9237 61446 9289 61498
rect 9301 61446 9353 61498
rect 9365 61446 9417 61498
rect 2320 61140 2372 61192
rect 1492 61047 1544 61056
rect 1492 61013 1501 61047
rect 1501 61013 1535 61047
rect 1535 61013 1544 61047
rect 1492 61004 1544 61013
rect 4213 60902 4265 60954
rect 4277 60902 4329 60954
rect 4341 60902 4393 60954
rect 4405 60902 4457 60954
rect 4469 60902 4521 60954
rect 7477 60902 7529 60954
rect 7541 60902 7593 60954
rect 7605 60902 7657 60954
rect 7669 60902 7721 60954
rect 7733 60902 7785 60954
rect 3240 60596 3292 60648
rect 10048 60571 10100 60580
rect 10048 60537 10057 60571
rect 10057 60537 10091 60571
rect 10091 60537 10100 60571
rect 10048 60528 10100 60537
rect 1400 60460 1452 60512
rect 2582 60358 2634 60410
rect 2646 60358 2698 60410
rect 2710 60358 2762 60410
rect 2774 60358 2826 60410
rect 2838 60358 2890 60410
rect 5845 60358 5897 60410
rect 5909 60358 5961 60410
rect 5973 60358 6025 60410
rect 6037 60358 6089 60410
rect 6101 60358 6153 60410
rect 9109 60358 9161 60410
rect 9173 60358 9225 60410
rect 9237 60358 9289 60410
rect 9301 60358 9353 60410
rect 9365 60358 9417 60410
rect 3424 60052 3476 60104
rect 9772 60052 9824 60104
rect 1492 59959 1544 59968
rect 1492 59925 1501 59959
rect 1501 59925 1535 59959
rect 1535 59925 1544 59959
rect 1492 59916 1544 59925
rect 10048 59959 10100 59968
rect 10048 59925 10057 59959
rect 10057 59925 10091 59959
rect 10091 59925 10100 59959
rect 10048 59916 10100 59925
rect 4213 59814 4265 59866
rect 4277 59814 4329 59866
rect 4341 59814 4393 59866
rect 4405 59814 4457 59866
rect 4469 59814 4521 59866
rect 7477 59814 7529 59866
rect 7541 59814 7593 59866
rect 7605 59814 7657 59866
rect 7669 59814 7721 59866
rect 7733 59814 7785 59866
rect 3608 59576 3660 59628
rect 9864 59619 9916 59628
rect 9864 59585 9873 59619
rect 9873 59585 9907 59619
rect 9907 59585 9916 59619
rect 9864 59576 9916 59585
rect 1400 59372 1452 59424
rect 10048 59415 10100 59424
rect 10048 59381 10057 59415
rect 10057 59381 10091 59415
rect 10091 59381 10100 59415
rect 10048 59372 10100 59381
rect 2582 59270 2634 59322
rect 2646 59270 2698 59322
rect 2710 59270 2762 59322
rect 2774 59270 2826 59322
rect 2838 59270 2890 59322
rect 5845 59270 5897 59322
rect 5909 59270 5961 59322
rect 5973 59270 6025 59322
rect 6037 59270 6089 59322
rect 6101 59270 6153 59322
rect 9109 59270 9161 59322
rect 9173 59270 9225 59322
rect 9237 59270 9289 59322
rect 9301 59270 9353 59322
rect 9365 59270 9417 59322
rect 1768 59100 1820 59152
rect 2136 59100 2188 59152
rect 1768 58964 1820 59016
rect 1492 58871 1544 58880
rect 1492 58837 1501 58871
rect 1501 58837 1535 58871
rect 1535 58837 1544 58871
rect 1492 58828 1544 58837
rect 4213 58726 4265 58778
rect 4277 58726 4329 58778
rect 4341 58726 4393 58778
rect 4405 58726 4457 58778
rect 4469 58726 4521 58778
rect 7477 58726 7529 58778
rect 7541 58726 7593 58778
rect 7605 58726 7657 58778
rect 7669 58726 7721 58778
rect 7733 58726 7785 58778
rect 1952 58488 2004 58540
rect 10048 58395 10100 58404
rect 10048 58361 10057 58395
rect 10057 58361 10091 58395
rect 10091 58361 10100 58395
rect 10048 58352 10100 58361
rect 1400 58284 1452 58336
rect 2582 58182 2634 58234
rect 2646 58182 2698 58234
rect 2710 58182 2762 58234
rect 2774 58182 2826 58234
rect 2838 58182 2890 58234
rect 5845 58182 5897 58234
rect 5909 58182 5961 58234
rect 5973 58182 6025 58234
rect 6037 58182 6089 58234
rect 6101 58182 6153 58234
rect 9109 58182 9161 58234
rect 9173 58182 9225 58234
rect 9237 58182 9289 58234
rect 9301 58182 9353 58234
rect 9365 58182 9417 58234
rect 1308 58012 1360 58064
rect 2228 58012 2280 58064
rect 1492 57876 1544 57928
rect 2228 57876 2280 57928
rect 2596 57876 2648 57928
rect 1492 57740 1544 57792
rect 8576 57808 8628 57860
rect 1952 57783 2004 57792
rect 1952 57749 1961 57783
rect 1961 57749 1995 57783
rect 1995 57749 2004 57783
rect 1952 57740 2004 57749
rect 2780 57740 2832 57792
rect 10048 57783 10100 57792
rect 10048 57749 10057 57783
rect 10057 57749 10091 57783
rect 10091 57749 10100 57783
rect 10048 57740 10100 57749
rect 4213 57638 4265 57690
rect 4277 57638 4329 57690
rect 4341 57638 4393 57690
rect 4405 57638 4457 57690
rect 4469 57638 4521 57690
rect 7477 57638 7529 57690
rect 7541 57638 7593 57690
rect 7605 57638 7657 57690
rect 7669 57638 7721 57690
rect 7733 57638 7785 57690
rect 1952 57536 2004 57588
rect 1676 57511 1728 57520
rect 1676 57477 1685 57511
rect 1685 57477 1719 57511
rect 1719 57477 1728 57511
rect 1676 57468 1728 57477
rect 3148 57468 3200 57520
rect 3332 57468 3384 57520
rect 1492 57400 1544 57452
rect 1952 57400 2004 57452
rect 2596 57400 2648 57452
rect 3516 57400 3568 57452
rect 7380 57332 7432 57384
rect 9864 57264 9916 57316
rect 2964 57196 3016 57248
rect 10048 57239 10100 57248
rect 10048 57205 10057 57239
rect 10057 57205 10091 57239
rect 10091 57205 10100 57239
rect 10048 57196 10100 57205
rect 2582 57094 2634 57146
rect 2646 57094 2698 57146
rect 2710 57094 2762 57146
rect 2774 57094 2826 57146
rect 2838 57094 2890 57146
rect 5845 57094 5897 57146
rect 5909 57094 5961 57146
rect 5973 57094 6025 57146
rect 6037 57094 6089 57146
rect 6101 57094 6153 57146
rect 9109 57094 9161 57146
rect 9173 57094 9225 57146
rect 9237 57094 9289 57146
rect 9301 57094 9353 57146
rect 9365 57094 9417 57146
rect 3240 56992 3292 57044
rect 3884 56992 3936 57044
rect 9772 56924 9824 56976
rect 1400 56831 1452 56840
rect 1400 56797 1409 56831
rect 1409 56797 1443 56831
rect 1443 56797 1452 56831
rect 1400 56788 1452 56797
rect 7288 56856 7340 56908
rect 1952 56788 2004 56840
rect 2688 56788 2740 56840
rect 3884 56788 3936 56840
rect 2044 56720 2096 56772
rect 3148 56720 3200 56772
rect 1860 56652 1912 56704
rect 1952 56652 2004 56704
rect 2228 56652 2280 56704
rect 2872 56652 2924 56704
rect 3976 56695 4028 56704
rect 3976 56661 3985 56695
rect 3985 56661 4019 56695
rect 4019 56661 4028 56695
rect 3976 56652 4028 56661
rect 4213 56550 4265 56602
rect 4277 56550 4329 56602
rect 4341 56550 4393 56602
rect 4405 56550 4457 56602
rect 4469 56550 4521 56602
rect 7477 56550 7529 56602
rect 7541 56550 7593 56602
rect 7605 56550 7657 56602
rect 7669 56550 7721 56602
rect 7733 56550 7785 56602
rect 1400 56355 1452 56364
rect 1400 56321 1409 56355
rect 1409 56321 1443 56355
rect 1443 56321 1452 56355
rect 1400 56312 1452 56321
rect 1676 56448 1728 56500
rect 2596 56448 2648 56500
rect 3608 56448 3660 56500
rect 4068 56448 4120 56500
rect 2688 56312 2740 56364
rect 2872 56244 2924 56296
rect 3056 56312 3108 56364
rect 3608 56312 3660 56364
rect 5816 56380 5868 56432
rect 3056 56176 3108 56228
rect 3976 56244 4028 56296
rect 8668 56176 8720 56228
rect 1860 56108 1912 56160
rect 10048 56151 10100 56160
rect 10048 56117 10057 56151
rect 10057 56117 10091 56151
rect 10091 56117 10100 56151
rect 10048 56108 10100 56117
rect 2582 56006 2634 56058
rect 2646 56006 2698 56058
rect 2710 56006 2762 56058
rect 2774 56006 2826 56058
rect 2838 56006 2890 56058
rect 5845 56006 5897 56058
rect 5909 56006 5961 56058
rect 5973 56006 6025 56058
rect 6037 56006 6089 56058
rect 6101 56006 6153 56058
rect 9109 56006 9161 56058
rect 9173 56006 9225 56058
rect 9237 56006 9289 56058
rect 9301 56006 9353 56058
rect 9365 56006 9417 56058
rect 1400 55768 1452 55820
rect 4068 55768 4120 55820
rect 2320 55700 2372 55752
rect 3056 55632 3108 55684
rect 3976 55607 4028 55616
rect 3976 55573 3985 55607
rect 3985 55573 4019 55607
rect 4019 55573 4028 55607
rect 3976 55564 4028 55573
rect 10048 55607 10100 55616
rect 10048 55573 10057 55607
rect 10057 55573 10091 55607
rect 10091 55573 10100 55607
rect 10048 55564 10100 55573
rect 4213 55462 4265 55514
rect 4277 55462 4329 55514
rect 4341 55462 4393 55514
rect 4405 55462 4457 55514
rect 4469 55462 4521 55514
rect 7477 55462 7529 55514
rect 7541 55462 7593 55514
rect 7605 55462 7657 55514
rect 7669 55462 7721 55514
rect 7733 55462 7785 55514
rect 2688 55360 2740 55412
rect 2964 55360 3016 55412
rect 1400 55267 1452 55276
rect 1400 55233 1409 55267
rect 1409 55233 1443 55267
rect 1443 55233 1452 55267
rect 1400 55224 1452 55233
rect 1676 55267 1728 55276
rect 1676 55233 1685 55267
rect 1685 55233 1719 55267
rect 1719 55233 1728 55267
rect 1676 55224 1728 55233
rect 1860 55224 1912 55276
rect 2044 55224 2096 55276
rect 8760 55224 8812 55276
rect 1584 55156 1636 55208
rect 4712 55156 4764 55208
rect 5540 55156 5592 55208
rect 1400 55088 1452 55140
rect 2688 55088 2740 55140
rect 2582 54918 2634 54970
rect 2646 54918 2698 54970
rect 2710 54918 2762 54970
rect 2774 54918 2826 54970
rect 2838 54918 2890 54970
rect 5845 54918 5897 54970
rect 5909 54918 5961 54970
rect 5973 54918 6025 54970
rect 6037 54918 6089 54970
rect 6101 54918 6153 54970
rect 9109 54918 9161 54970
rect 9173 54918 9225 54970
rect 9237 54918 9289 54970
rect 9301 54918 9353 54970
rect 9365 54918 9417 54970
rect 1400 54612 1452 54664
rect 10140 54655 10192 54664
rect 10140 54621 10149 54655
rect 10149 54621 10183 54655
rect 10183 54621 10192 54655
rect 10140 54612 10192 54621
rect 1492 54519 1544 54528
rect 1492 54485 1501 54519
rect 1501 54485 1535 54519
rect 1535 54485 1544 54519
rect 1492 54476 1544 54485
rect 9956 54519 10008 54528
rect 9956 54485 9965 54519
rect 9965 54485 9999 54519
rect 9999 54485 10008 54519
rect 9956 54476 10008 54485
rect 4213 54374 4265 54426
rect 4277 54374 4329 54426
rect 4341 54374 4393 54426
rect 4405 54374 4457 54426
rect 4469 54374 4521 54426
rect 7477 54374 7529 54426
rect 7541 54374 7593 54426
rect 7605 54374 7657 54426
rect 7669 54374 7721 54426
rect 7733 54374 7785 54426
rect 3148 54204 3200 54256
rect 3240 54136 3292 54188
rect 3976 54179 4028 54188
rect 3976 54145 3985 54179
rect 3985 54145 4019 54179
rect 4019 54145 4028 54179
rect 3976 54136 4028 54145
rect 10140 54179 10192 54188
rect 10140 54145 10149 54179
rect 10149 54145 10183 54179
rect 10183 54145 10192 54179
rect 10140 54136 10192 54145
rect 2964 54068 3016 54120
rect 3148 54068 3200 54120
rect 3516 54068 3568 54120
rect 1492 53975 1544 53984
rect 1492 53941 1501 53975
rect 1501 53941 1535 53975
rect 1535 53941 1544 53975
rect 1492 53932 1544 53941
rect 9864 53932 9916 53984
rect 2582 53830 2634 53882
rect 2646 53830 2698 53882
rect 2710 53830 2762 53882
rect 2774 53830 2826 53882
rect 2838 53830 2890 53882
rect 5845 53830 5897 53882
rect 5909 53830 5961 53882
rect 5973 53830 6025 53882
rect 6037 53830 6089 53882
rect 6101 53830 6153 53882
rect 9109 53830 9161 53882
rect 9173 53830 9225 53882
rect 9237 53830 9289 53882
rect 9301 53830 9353 53882
rect 9365 53830 9417 53882
rect 3056 53592 3108 53644
rect 2228 53524 2280 53576
rect 9956 53524 10008 53576
rect 10140 53567 10192 53576
rect 10140 53533 10149 53567
rect 10149 53533 10183 53567
rect 10183 53533 10192 53567
rect 10140 53524 10192 53533
rect 3056 53388 3108 53440
rect 9956 53431 10008 53440
rect 9956 53397 9965 53431
rect 9965 53397 9999 53431
rect 9999 53397 10008 53431
rect 9956 53388 10008 53397
rect 4213 53286 4265 53338
rect 4277 53286 4329 53338
rect 4341 53286 4393 53338
rect 4405 53286 4457 53338
rect 4469 53286 4521 53338
rect 7477 53286 7529 53338
rect 7541 53286 7593 53338
rect 7605 53286 7657 53338
rect 7669 53286 7721 53338
rect 7733 53286 7785 53338
rect 1492 53184 1544 53236
rect 3792 53184 3844 53236
rect 848 53116 900 53168
rect 1952 53048 2004 53100
rect 2780 53048 2832 53100
rect 3056 53091 3108 53100
rect 3056 53057 3065 53091
rect 3065 53057 3099 53091
rect 3099 53057 3108 53091
rect 3056 53048 3108 53057
rect 9864 53048 9916 53100
rect 3516 52980 3568 53032
rect 204 52912 256 52964
rect 1492 52887 1544 52896
rect 1492 52853 1501 52887
rect 1501 52853 1535 52887
rect 1535 52853 1544 52887
rect 1492 52844 1544 52853
rect 3240 52844 3292 52896
rect 2582 52742 2634 52794
rect 2646 52742 2698 52794
rect 2710 52742 2762 52794
rect 2774 52742 2826 52794
rect 2838 52742 2890 52794
rect 5845 52742 5897 52794
rect 5909 52742 5961 52794
rect 5973 52742 6025 52794
rect 6037 52742 6089 52794
rect 6101 52742 6153 52794
rect 9109 52742 9161 52794
rect 9173 52742 9225 52794
rect 9237 52742 9289 52794
rect 9301 52742 9353 52794
rect 9365 52742 9417 52794
rect 1308 52640 1360 52692
rect 1676 52640 1728 52692
rect 2412 52683 2464 52692
rect 2412 52649 2421 52683
rect 2421 52649 2455 52683
rect 2455 52649 2464 52683
rect 2412 52640 2464 52649
rect 3700 52640 3752 52692
rect 756 52572 808 52624
rect 3148 52504 3200 52556
rect 1492 52343 1544 52352
rect 1492 52309 1501 52343
rect 1501 52309 1535 52343
rect 1535 52309 1544 52343
rect 1492 52300 1544 52309
rect 3240 52479 3292 52488
rect 3240 52445 3249 52479
rect 3249 52445 3283 52479
rect 3283 52445 3292 52479
rect 3240 52436 3292 52445
rect 9956 52436 10008 52488
rect 10140 52479 10192 52488
rect 10140 52445 10149 52479
rect 10149 52445 10183 52479
rect 10183 52445 10192 52479
rect 10140 52436 10192 52445
rect 5448 52368 5500 52420
rect 3148 52300 3200 52352
rect 3608 52300 3660 52352
rect 4068 52300 4120 52352
rect 9496 52300 9548 52352
rect 4213 52198 4265 52250
rect 4277 52198 4329 52250
rect 4341 52198 4393 52250
rect 4405 52198 4457 52250
rect 4469 52198 4521 52250
rect 7477 52198 7529 52250
rect 7541 52198 7593 52250
rect 7605 52198 7657 52250
rect 7669 52198 7721 52250
rect 7733 52198 7785 52250
rect 2136 52096 2188 52148
rect 3424 52096 3476 52148
rect 8024 52028 8076 52080
rect 2136 51960 2188 52012
rect 2504 51960 2556 52012
rect 4068 51960 4120 52012
rect 10140 52003 10192 52012
rect 10140 51969 10149 52003
rect 10149 51969 10183 52003
rect 10183 51969 10192 52003
rect 10140 51960 10192 51969
rect 3424 51892 3476 51944
rect 2228 51756 2280 51808
rect 2780 51824 2832 51876
rect 9956 51799 10008 51808
rect 9956 51765 9965 51799
rect 9965 51765 9999 51799
rect 9999 51765 10008 51799
rect 9956 51756 10008 51765
rect 2582 51654 2634 51706
rect 2646 51654 2698 51706
rect 2710 51654 2762 51706
rect 2774 51654 2826 51706
rect 2838 51654 2890 51706
rect 5845 51654 5897 51706
rect 5909 51654 5961 51706
rect 5973 51654 6025 51706
rect 6037 51654 6089 51706
rect 6101 51654 6153 51706
rect 9109 51654 9161 51706
rect 9173 51654 9225 51706
rect 9237 51654 9289 51706
rect 9301 51654 9353 51706
rect 9365 51654 9417 51706
rect 2412 51552 2464 51604
rect 2596 51484 2648 51536
rect 1676 51391 1728 51400
rect 1676 51357 1685 51391
rect 1685 51357 1719 51391
rect 1719 51357 1728 51391
rect 2136 51416 2188 51468
rect 2320 51416 2372 51468
rect 1676 51348 1728 51357
rect 2228 51348 2280 51400
rect 2412 51391 2464 51400
rect 2412 51357 2421 51391
rect 2421 51357 2455 51391
rect 2455 51357 2464 51391
rect 2412 51348 2464 51357
rect 5816 51416 5868 51468
rect 2964 51348 3016 51400
rect 3240 51348 3292 51400
rect 9496 51348 9548 51400
rect 1492 51212 1544 51264
rect 1584 51212 1636 51264
rect 2136 51212 2188 51264
rect 3240 51212 3292 51264
rect 4896 51212 4948 51264
rect 4213 51110 4265 51162
rect 4277 51110 4329 51162
rect 4341 51110 4393 51162
rect 4405 51110 4457 51162
rect 4469 51110 4521 51162
rect 7477 51110 7529 51162
rect 7541 51110 7593 51162
rect 7605 51110 7657 51162
rect 7669 51110 7721 51162
rect 7733 51110 7785 51162
rect 2412 51008 2464 51060
rect 3608 51008 3660 51060
rect 1676 50983 1728 50992
rect 1676 50949 1685 50983
rect 1685 50949 1719 50983
rect 1719 50949 1728 50983
rect 1676 50940 1728 50949
rect 1400 50915 1452 50924
rect 1400 50881 1409 50915
rect 1409 50881 1443 50915
rect 1443 50881 1452 50915
rect 1400 50872 1452 50881
rect 2320 50940 2372 50992
rect 2412 50915 2464 50924
rect 2412 50881 2421 50915
rect 2421 50881 2455 50915
rect 2455 50881 2464 50915
rect 2412 50872 2464 50881
rect 3056 50804 3108 50856
rect 3976 50872 4028 50924
rect 9956 51008 10008 51060
rect 4896 50915 4948 50924
rect 4896 50881 4905 50915
rect 4905 50881 4939 50915
rect 4939 50881 4948 50915
rect 4896 50872 4948 50881
rect 10140 50915 10192 50924
rect 10140 50881 10149 50915
rect 10149 50881 10183 50915
rect 10183 50881 10192 50915
rect 10140 50872 10192 50881
rect 2780 50736 2832 50788
rect 3332 50736 3384 50788
rect 4068 50711 4120 50720
rect 4068 50677 4077 50711
rect 4077 50677 4111 50711
rect 4111 50677 4120 50711
rect 4068 50668 4120 50677
rect 4160 50668 4212 50720
rect 9956 50711 10008 50720
rect 9956 50677 9965 50711
rect 9965 50677 9999 50711
rect 9999 50677 10008 50711
rect 9956 50668 10008 50677
rect 2582 50566 2634 50618
rect 2646 50566 2698 50618
rect 2710 50566 2762 50618
rect 2774 50566 2826 50618
rect 2838 50566 2890 50618
rect 5845 50566 5897 50618
rect 5909 50566 5961 50618
rect 5973 50566 6025 50618
rect 6037 50566 6089 50618
rect 6101 50566 6153 50618
rect 9109 50566 9161 50618
rect 9173 50566 9225 50618
rect 9237 50566 9289 50618
rect 9301 50566 9353 50618
rect 9365 50566 9417 50618
rect 3056 50464 3108 50516
rect 8116 50464 8168 50516
rect 3424 50328 3476 50380
rect 4160 50328 4212 50380
rect 1400 50303 1452 50312
rect 1400 50269 1409 50303
rect 1409 50269 1443 50303
rect 1443 50269 1452 50303
rect 1400 50260 1452 50269
rect 1492 50260 1544 50312
rect 2320 50260 2372 50312
rect 3056 50260 3108 50312
rect 9956 50260 10008 50312
rect 10140 50303 10192 50312
rect 10140 50269 10149 50303
rect 10149 50269 10183 50303
rect 10183 50269 10192 50303
rect 10140 50260 10192 50269
rect 3424 50192 3476 50244
rect 2504 50167 2556 50176
rect 2504 50133 2513 50167
rect 2513 50133 2547 50167
rect 2547 50133 2556 50167
rect 2504 50124 2556 50133
rect 3976 50124 4028 50176
rect 6276 50124 6328 50176
rect 9956 50167 10008 50176
rect 9956 50133 9965 50167
rect 9965 50133 9999 50167
rect 9999 50133 10008 50167
rect 9956 50124 10008 50133
rect 4213 50022 4265 50074
rect 4277 50022 4329 50074
rect 4341 50022 4393 50074
rect 4405 50022 4457 50074
rect 4469 50022 4521 50074
rect 7477 50022 7529 50074
rect 7541 50022 7593 50074
rect 7605 50022 7657 50074
rect 7669 50022 7721 50074
rect 7733 50022 7785 50074
rect 1768 49920 1820 49972
rect 1768 49784 1820 49836
rect 4712 49920 4764 49972
rect 1492 49691 1544 49700
rect 1492 49657 1501 49691
rect 1501 49657 1535 49691
rect 1535 49657 1544 49691
rect 1492 49648 1544 49657
rect 3516 49784 3568 49836
rect 3976 49784 4028 49836
rect 9956 49784 10008 49836
rect 4068 49716 4120 49768
rect 4988 49716 5040 49768
rect 3332 49648 3384 49700
rect 5448 49648 5500 49700
rect 10140 49648 10192 49700
rect 4252 49580 4304 49632
rect 2582 49478 2634 49530
rect 2646 49478 2698 49530
rect 2710 49478 2762 49530
rect 2774 49478 2826 49530
rect 2838 49478 2890 49530
rect 5845 49478 5897 49530
rect 5909 49478 5961 49530
rect 5973 49478 6025 49530
rect 6037 49478 6089 49530
rect 6101 49478 6153 49530
rect 9109 49478 9161 49530
rect 9173 49478 9225 49530
rect 9237 49478 9289 49530
rect 9301 49478 9353 49530
rect 9365 49478 9417 49530
rect 1860 49376 1912 49428
rect 664 49240 716 49292
rect 1860 49172 1912 49224
rect 4252 49215 4304 49224
rect 4252 49181 4261 49215
rect 4261 49181 4295 49215
rect 4295 49181 4304 49215
rect 4252 49172 4304 49181
rect 3332 49104 3384 49156
rect 1492 49079 1544 49088
rect 1492 49045 1501 49079
rect 1501 49045 1535 49079
rect 1535 49045 1544 49079
rect 1492 49036 1544 49045
rect 4213 48934 4265 48986
rect 4277 48934 4329 48986
rect 4341 48934 4393 48986
rect 4405 48934 4457 48986
rect 4469 48934 4521 48986
rect 7477 48934 7529 48986
rect 7541 48934 7593 48986
rect 7605 48934 7657 48986
rect 7669 48934 7721 48986
rect 7733 48934 7785 48986
rect 3792 48875 3844 48884
rect 3792 48841 3801 48875
rect 3801 48841 3835 48875
rect 3835 48841 3844 48875
rect 3792 48832 3844 48841
rect 3516 48696 3568 48748
rect 10140 48739 10192 48748
rect 572 48628 624 48680
rect 10140 48705 10149 48739
rect 10149 48705 10183 48739
rect 10183 48705 10192 48739
rect 10140 48696 10192 48705
rect 1492 48603 1544 48612
rect 1492 48569 1501 48603
rect 1501 48569 1535 48603
rect 1535 48569 1544 48603
rect 1492 48560 1544 48569
rect 3792 48492 3844 48544
rect 9956 48535 10008 48544
rect 9956 48501 9965 48535
rect 9965 48501 9999 48535
rect 9999 48501 10008 48535
rect 9956 48492 10008 48501
rect 2582 48390 2634 48442
rect 2646 48390 2698 48442
rect 2710 48390 2762 48442
rect 2774 48390 2826 48442
rect 2838 48390 2890 48442
rect 5845 48390 5897 48442
rect 5909 48390 5961 48442
rect 5973 48390 6025 48442
rect 6037 48390 6089 48442
rect 6101 48390 6153 48442
rect 9109 48390 9161 48442
rect 9173 48390 9225 48442
rect 9237 48390 9289 48442
rect 9301 48390 9353 48442
rect 9365 48390 9417 48442
rect 2320 48084 2372 48136
rect 10140 48127 10192 48136
rect 10140 48093 10149 48127
rect 10149 48093 10183 48127
rect 10183 48093 10192 48127
rect 10140 48084 10192 48093
rect 1492 47991 1544 48000
rect 1492 47957 1501 47991
rect 1501 47957 1535 47991
rect 1535 47957 1544 47991
rect 1492 47948 1544 47957
rect 9864 47948 9916 48000
rect 4213 47846 4265 47898
rect 4277 47846 4329 47898
rect 4341 47846 4393 47898
rect 4405 47846 4457 47898
rect 4469 47846 4521 47898
rect 7477 47846 7529 47898
rect 7541 47846 7593 47898
rect 7605 47846 7657 47898
rect 7669 47846 7721 47898
rect 7733 47846 7785 47898
rect 756 47608 808 47660
rect 1676 47651 1728 47660
rect 1676 47617 1685 47651
rect 1685 47617 1719 47651
rect 1719 47617 1728 47651
rect 1676 47608 1728 47617
rect 3332 47651 3384 47660
rect 3332 47617 3341 47651
rect 3341 47617 3375 47651
rect 3375 47617 3384 47651
rect 3332 47608 3384 47617
rect 9956 47608 10008 47660
rect 3608 47583 3660 47592
rect 3608 47549 3617 47583
rect 3617 47549 3651 47583
rect 3651 47549 3660 47583
rect 3608 47540 3660 47549
rect 1492 47515 1544 47524
rect 1492 47481 1501 47515
rect 1501 47481 1535 47515
rect 1535 47481 1544 47515
rect 1492 47472 1544 47481
rect 848 47404 900 47456
rect 4160 47447 4212 47456
rect 4160 47413 4169 47447
rect 4169 47413 4203 47447
rect 4203 47413 4212 47447
rect 4160 47404 4212 47413
rect 2582 47302 2634 47354
rect 2646 47302 2698 47354
rect 2710 47302 2762 47354
rect 2774 47302 2826 47354
rect 2838 47302 2890 47354
rect 5845 47302 5897 47354
rect 5909 47302 5961 47354
rect 5973 47302 6025 47354
rect 6037 47302 6089 47354
rect 6101 47302 6153 47354
rect 9109 47302 9161 47354
rect 9173 47302 9225 47354
rect 9237 47302 9289 47354
rect 9301 47302 9353 47354
rect 9365 47302 9417 47354
rect 1492 47175 1544 47184
rect 1492 47141 1501 47175
rect 1501 47141 1535 47175
rect 1535 47141 1544 47175
rect 1492 47132 1544 47141
rect 3332 46996 3384 47048
rect 10140 47039 10192 47048
rect 10140 47005 10149 47039
rect 10149 47005 10183 47039
rect 10183 47005 10192 47039
rect 10140 46996 10192 47005
rect 4068 46860 4120 46912
rect 4213 46758 4265 46810
rect 4277 46758 4329 46810
rect 4341 46758 4393 46810
rect 4405 46758 4457 46810
rect 4469 46758 4521 46810
rect 7477 46758 7529 46810
rect 7541 46758 7593 46810
rect 7605 46758 7657 46810
rect 7669 46758 7721 46810
rect 7733 46758 7785 46810
rect 2136 46656 2188 46708
rect 1584 46520 1636 46572
rect 2136 46563 2188 46572
rect 2136 46529 2145 46563
rect 2145 46529 2179 46563
rect 2179 46529 2188 46563
rect 2136 46520 2188 46529
rect 3976 46588 4028 46640
rect 112 46452 164 46504
rect 9864 46520 9916 46572
rect 10140 46563 10192 46572
rect 10140 46529 10149 46563
rect 10149 46529 10183 46563
rect 10183 46529 10192 46563
rect 10140 46520 10192 46529
rect 3976 46384 4028 46436
rect 7932 46384 7984 46436
rect 1492 46359 1544 46368
rect 1492 46325 1501 46359
rect 1501 46325 1535 46359
rect 1535 46325 1544 46359
rect 1492 46316 1544 46325
rect 7104 46316 7156 46368
rect 7380 46316 7432 46368
rect 9956 46359 10008 46368
rect 9956 46325 9965 46359
rect 9965 46325 9999 46359
rect 9999 46325 10008 46359
rect 9956 46316 10008 46325
rect 2582 46214 2634 46266
rect 2646 46214 2698 46266
rect 2710 46214 2762 46266
rect 2774 46214 2826 46266
rect 2838 46214 2890 46266
rect 5845 46214 5897 46266
rect 5909 46214 5961 46266
rect 5973 46214 6025 46266
rect 6037 46214 6089 46266
rect 6101 46214 6153 46266
rect 9109 46214 9161 46266
rect 9173 46214 9225 46266
rect 9237 46214 9289 46266
rect 9301 46214 9353 46266
rect 9365 46214 9417 46266
rect 2228 46112 2280 46164
rect 3884 46112 3936 46164
rect 3516 46044 3568 46096
rect 3700 46044 3752 46096
rect 7840 46044 7892 46096
rect 8116 46044 8168 46096
rect 2136 45951 2188 45960
rect 2136 45917 2145 45951
rect 2145 45917 2179 45951
rect 2179 45917 2188 45951
rect 2136 45908 2188 45917
rect 2228 45840 2280 45892
rect 1492 45815 1544 45824
rect 1492 45781 1501 45815
rect 1501 45781 1535 45815
rect 1535 45781 1544 45815
rect 1492 45772 1544 45781
rect 3976 45976 4028 46028
rect 2596 45840 2648 45892
rect 3056 45908 3108 45960
rect 3516 45908 3568 45960
rect 4068 45951 4120 45960
rect 4068 45917 4077 45951
rect 4077 45917 4111 45951
rect 4111 45917 4120 45951
rect 4068 45908 4120 45917
rect 10140 45951 10192 45960
rect 10140 45917 10149 45951
rect 10149 45917 10183 45951
rect 10183 45917 10192 45951
rect 10140 45908 10192 45917
rect 3792 45883 3844 45892
rect 3792 45849 3801 45883
rect 3801 45849 3835 45883
rect 3835 45849 3844 45883
rect 3792 45840 3844 45849
rect 3976 45772 4028 45824
rect 9864 45772 9916 45824
rect 4213 45670 4265 45722
rect 4277 45670 4329 45722
rect 4341 45670 4393 45722
rect 4405 45670 4457 45722
rect 4469 45670 4521 45722
rect 7477 45670 7529 45722
rect 7541 45670 7593 45722
rect 7605 45670 7657 45722
rect 7669 45670 7721 45722
rect 7733 45670 7785 45722
rect 2504 45500 2556 45552
rect 1400 45432 1452 45484
rect 2596 45432 2648 45484
rect 9956 45432 10008 45484
rect 2688 45407 2740 45416
rect 2688 45373 2697 45407
rect 2697 45373 2731 45407
rect 2731 45373 2740 45407
rect 2688 45364 2740 45373
rect 4068 45364 4120 45416
rect 1492 45271 1544 45280
rect 1492 45237 1501 45271
rect 1501 45237 1535 45271
rect 1535 45237 1544 45271
rect 1492 45228 1544 45237
rect 3976 45228 4028 45280
rect 6736 45228 6788 45280
rect 2582 45126 2634 45178
rect 2646 45126 2698 45178
rect 2710 45126 2762 45178
rect 2774 45126 2826 45178
rect 2838 45126 2890 45178
rect 5845 45126 5897 45178
rect 5909 45126 5961 45178
rect 5973 45126 6025 45178
rect 6037 45126 6089 45178
rect 6101 45126 6153 45178
rect 9109 45126 9161 45178
rect 9173 45126 9225 45178
rect 9237 45126 9289 45178
rect 9301 45126 9353 45178
rect 9365 45126 9417 45178
rect 2044 45024 2096 45076
rect 2964 45024 3016 45076
rect 20 44956 72 45008
rect 2136 44863 2188 44872
rect 2136 44829 2145 44863
rect 2145 44829 2179 44863
rect 2179 44829 2188 44863
rect 2136 44820 2188 44829
rect 2504 44888 2556 44940
rect 3792 44820 3844 44872
rect 1492 44727 1544 44736
rect 1492 44693 1501 44727
rect 1501 44693 1535 44727
rect 1535 44693 1544 44727
rect 1492 44684 1544 44693
rect 1860 44684 1912 44736
rect 2136 44684 2188 44736
rect 9864 44820 9916 44872
rect 10140 44863 10192 44872
rect 10140 44829 10149 44863
rect 10149 44829 10183 44863
rect 10183 44829 10192 44863
rect 10140 44820 10192 44829
rect 6368 44752 6420 44804
rect 2780 44684 2832 44736
rect 3516 44684 3568 44736
rect 3792 44684 3844 44736
rect 9956 44727 10008 44736
rect 9956 44693 9965 44727
rect 9965 44693 9999 44727
rect 9999 44693 10008 44727
rect 9956 44684 10008 44693
rect 4213 44582 4265 44634
rect 4277 44582 4329 44634
rect 4341 44582 4393 44634
rect 4405 44582 4457 44634
rect 4469 44582 4521 44634
rect 7477 44582 7529 44634
rect 7541 44582 7593 44634
rect 7605 44582 7657 44634
rect 7669 44582 7721 44634
rect 7733 44582 7785 44634
rect 10140 44387 10192 44396
rect 10140 44353 10149 44387
rect 10149 44353 10183 44387
rect 10183 44353 10192 44387
rect 10140 44344 10192 44353
rect 2044 44276 2096 44328
rect 1492 44183 1544 44192
rect 1492 44149 1501 44183
rect 1501 44149 1535 44183
rect 1535 44149 1544 44183
rect 1492 44140 1544 44149
rect 9864 44140 9916 44192
rect 2582 44038 2634 44090
rect 2646 44038 2698 44090
rect 2710 44038 2762 44090
rect 2774 44038 2826 44090
rect 2838 44038 2890 44090
rect 5845 44038 5897 44090
rect 5909 44038 5961 44090
rect 5973 44038 6025 44090
rect 6037 44038 6089 44090
rect 6101 44038 6153 44090
rect 9109 44038 9161 44090
rect 9173 44038 9225 44090
rect 9237 44038 9289 44090
rect 9301 44038 9353 44090
rect 9365 44038 9417 44090
rect 2504 43732 2556 43784
rect 10140 43775 10192 43784
rect 10140 43741 10149 43775
rect 10149 43741 10183 43775
rect 10183 43741 10192 43775
rect 10140 43732 10192 43741
rect 1492 43639 1544 43648
rect 1492 43605 1501 43639
rect 1501 43605 1535 43639
rect 1535 43605 1544 43639
rect 1492 43596 1544 43605
rect 9772 43596 9824 43648
rect 4213 43494 4265 43546
rect 4277 43494 4329 43546
rect 4341 43494 4393 43546
rect 4405 43494 4457 43546
rect 4469 43494 4521 43546
rect 7477 43494 7529 43546
rect 7541 43494 7593 43546
rect 7605 43494 7657 43546
rect 7669 43494 7721 43546
rect 7733 43494 7785 43546
rect 3332 43256 3384 43308
rect 9956 43256 10008 43308
rect 1492 43095 1544 43104
rect 1492 43061 1501 43095
rect 1501 43061 1535 43095
rect 1535 43061 1544 43095
rect 1492 43052 1544 43061
rect 3516 43052 3568 43104
rect 2582 42950 2634 43002
rect 2646 42950 2698 43002
rect 2710 42950 2762 43002
rect 2774 42950 2826 43002
rect 2838 42950 2890 43002
rect 5845 42950 5897 43002
rect 5909 42950 5961 43002
rect 5973 42950 6025 43002
rect 6037 42950 6089 43002
rect 6101 42950 6153 43002
rect 9109 42950 9161 43002
rect 9173 42950 9225 43002
rect 9237 42950 9289 43002
rect 9301 42950 9353 43002
rect 9365 42950 9417 43002
rect 4068 42755 4120 42764
rect 4068 42721 4077 42755
rect 4077 42721 4111 42755
rect 4111 42721 4120 42755
rect 4068 42712 4120 42721
rect 1860 42644 1912 42696
rect 3976 42644 4028 42696
rect 9496 42644 9548 42696
rect 10140 42687 10192 42696
rect 10140 42653 10149 42687
rect 10149 42653 10183 42687
rect 10183 42653 10192 42687
rect 10140 42644 10192 42653
rect 1492 42551 1544 42560
rect 1492 42517 1501 42551
rect 1501 42517 1535 42551
rect 1535 42517 1544 42551
rect 1492 42508 1544 42517
rect 9956 42551 10008 42560
rect 9956 42517 9965 42551
rect 9965 42517 9999 42551
rect 9999 42517 10008 42551
rect 9956 42508 10008 42517
rect 4213 42406 4265 42458
rect 4277 42406 4329 42458
rect 4341 42406 4393 42458
rect 4405 42406 4457 42458
rect 4469 42406 4521 42458
rect 7477 42406 7529 42458
rect 7541 42406 7593 42458
rect 7605 42406 7657 42458
rect 7669 42406 7721 42458
rect 7733 42406 7785 42458
rect 1400 42304 1452 42356
rect 1400 42168 1452 42220
rect 9864 42168 9916 42220
rect 10140 42211 10192 42220
rect 10140 42177 10149 42211
rect 10149 42177 10183 42211
rect 10183 42177 10192 42211
rect 10140 42168 10192 42177
rect 1492 42007 1544 42016
rect 1492 41973 1501 42007
rect 1501 41973 1535 42007
rect 1535 41973 1544 42007
rect 1492 41964 1544 41973
rect 3976 42007 4028 42016
rect 3976 41973 3985 42007
rect 3985 41973 4019 42007
rect 4019 41973 4028 42007
rect 3976 41964 4028 41973
rect 9864 41964 9916 42016
rect 2582 41862 2634 41914
rect 2646 41862 2698 41914
rect 2710 41862 2762 41914
rect 2774 41862 2826 41914
rect 2838 41862 2890 41914
rect 5845 41862 5897 41914
rect 5909 41862 5961 41914
rect 5973 41862 6025 41914
rect 6037 41862 6089 41914
rect 6101 41862 6153 41914
rect 9109 41862 9161 41914
rect 9173 41862 9225 41914
rect 9237 41862 9289 41914
rect 9301 41862 9353 41914
rect 9365 41862 9417 41914
rect 1308 41760 1360 41812
rect 4068 41692 4120 41744
rect 2136 41599 2188 41608
rect 2136 41565 2145 41599
rect 2145 41565 2179 41599
rect 2179 41565 2188 41599
rect 2136 41556 2188 41565
rect 2780 41556 2832 41608
rect 3516 41556 3568 41608
rect 9772 41556 9824 41608
rect 1308 41488 1360 41540
rect 2688 41488 2740 41540
rect 4160 41488 4212 41540
rect 1492 41463 1544 41472
rect 1492 41429 1501 41463
rect 1501 41429 1535 41463
rect 1535 41429 1544 41463
rect 1492 41420 1544 41429
rect 4213 41318 4265 41370
rect 4277 41318 4329 41370
rect 4341 41318 4393 41370
rect 4405 41318 4457 41370
rect 4469 41318 4521 41370
rect 7477 41318 7529 41370
rect 7541 41318 7593 41370
rect 7605 41318 7657 41370
rect 7669 41318 7721 41370
rect 7733 41318 7785 41370
rect 1308 41216 1360 41268
rect 1492 41216 1544 41268
rect 1952 41216 2004 41268
rect 3148 41216 3200 41268
rect 3516 41216 3568 41268
rect 2136 41123 2188 41132
rect 2136 41089 2145 41123
rect 2145 41089 2179 41123
rect 2179 41089 2188 41123
rect 2136 41080 2188 41089
rect 2688 41080 2740 41132
rect 3884 41148 3936 41200
rect 6460 41148 6512 41200
rect 6644 41148 6696 41200
rect 3976 41080 4028 41132
rect 9956 41080 10008 41132
rect 10140 41123 10192 41132
rect 10140 41089 10149 41123
rect 10149 41089 10183 41123
rect 10183 41089 10192 41123
rect 10140 41080 10192 41089
rect 1492 40919 1544 40928
rect 1492 40885 1501 40919
rect 1501 40885 1535 40919
rect 1535 40885 1544 40919
rect 1492 40876 1544 40885
rect 3884 40944 3936 40996
rect 4436 40876 4488 40928
rect 6552 40876 6604 40928
rect 9956 40919 10008 40928
rect 9956 40885 9965 40919
rect 9965 40885 9999 40919
rect 9999 40885 10008 40919
rect 9956 40876 10008 40885
rect 2582 40774 2634 40826
rect 2646 40774 2698 40826
rect 2710 40774 2762 40826
rect 2774 40774 2826 40826
rect 2838 40774 2890 40826
rect 5845 40774 5897 40826
rect 5909 40774 5961 40826
rect 5973 40774 6025 40826
rect 6037 40774 6089 40826
rect 6101 40774 6153 40826
rect 9109 40774 9161 40826
rect 9173 40774 9225 40826
rect 9237 40774 9289 40826
rect 9301 40774 9353 40826
rect 9365 40774 9417 40826
rect 1400 40672 1452 40724
rect 3608 40672 3660 40724
rect 4436 40672 4488 40724
rect 1584 40468 1636 40520
rect 2136 40511 2188 40520
rect 2136 40477 2145 40511
rect 2145 40477 2179 40511
rect 2179 40477 2188 40511
rect 2136 40468 2188 40477
rect 2872 40468 2924 40520
rect 1492 40375 1544 40384
rect 1492 40341 1501 40375
rect 1501 40341 1535 40375
rect 1535 40341 1544 40375
rect 1492 40332 1544 40341
rect 4620 40604 4672 40656
rect 5172 40604 5224 40656
rect 5080 40536 5132 40588
rect 5356 40536 5408 40588
rect 9864 40468 9916 40520
rect 10140 40511 10192 40520
rect 10140 40477 10149 40511
rect 10149 40477 10183 40511
rect 10183 40477 10192 40511
rect 10140 40468 10192 40477
rect 6828 40332 6880 40384
rect 9864 40332 9916 40384
rect 4213 40230 4265 40282
rect 4277 40230 4329 40282
rect 4341 40230 4393 40282
rect 4405 40230 4457 40282
rect 4469 40230 4521 40282
rect 7477 40230 7529 40282
rect 7541 40230 7593 40282
rect 7605 40230 7657 40282
rect 7669 40230 7721 40282
rect 7733 40230 7785 40282
rect 3976 40128 4028 40180
rect 5356 40128 5408 40180
rect 1400 40035 1452 40044
rect 1400 40001 1409 40035
rect 1409 40001 1443 40035
rect 1443 40001 1452 40035
rect 1400 39992 1452 40001
rect 2596 40035 2648 40044
rect 2596 40001 2605 40035
rect 2605 40001 2639 40035
rect 2639 40001 2648 40035
rect 2596 39992 2648 40001
rect 2872 40035 2924 40044
rect 2872 40001 2881 40035
rect 2881 40001 2915 40035
rect 2915 40001 2924 40035
rect 2872 39992 2924 40001
rect 9956 40060 10008 40112
rect 10140 40035 10192 40044
rect 10140 40001 10149 40035
rect 10149 40001 10183 40035
rect 10183 40001 10192 40035
rect 10140 39992 10192 40001
rect 5540 39856 5592 39908
rect 5080 39788 5132 39840
rect 9956 39831 10008 39840
rect 9956 39797 9965 39831
rect 9965 39797 9999 39831
rect 9999 39797 10008 39831
rect 9956 39788 10008 39797
rect 2582 39686 2634 39738
rect 2646 39686 2698 39738
rect 2710 39686 2762 39738
rect 2774 39686 2826 39738
rect 2838 39686 2890 39738
rect 5845 39686 5897 39738
rect 5909 39686 5961 39738
rect 5973 39686 6025 39738
rect 6037 39686 6089 39738
rect 6101 39686 6153 39738
rect 9109 39686 9161 39738
rect 9173 39686 9225 39738
rect 9237 39686 9289 39738
rect 9301 39686 9353 39738
rect 9365 39686 9417 39738
rect 2412 39584 2464 39636
rect 5264 39516 5316 39568
rect 2412 39448 2464 39500
rect 1400 39423 1452 39432
rect 1400 39389 1409 39423
rect 1409 39389 1443 39423
rect 1443 39389 1452 39423
rect 1400 39380 1452 39389
rect 2136 39423 2188 39432
rect 2136 39389 2145 39423
rect 2145 39389 2179 39423
rect 2179 39389 2188 39423
rect 2136 39380 2188 39389
rect 296 39312 348 39364
rect 9864 39380 9916 39432
rect 4213 39142 4265 39194
rect 4277 39142 4329 39194
rect 4341 39142 4393 39194
rect 4405 39142 4457 39194
rect 4469 39142 4521 39194
rect 7477 39142 7529 39194
rect 7541 39142 7593 39194
rect 7605 39142 7657 39194
rect 7669 39142 7721 39194
rect 7733 39142 7785 39194
rect 1124 39040 1176 39092
rect 1768 39040 1820 39092
rect 3148 39040 3200 39092
rect 1400 38947 1452 38956
rect 1400 38913 1409 38947
rect 1409 38913 1443 38947
rect 1443 38913 1452 38947
rect 1400 38904 1452 38913
rect 2136 38947 2188 38956
rect 2136 38913 2145 38947
rect 2145 38913 2179 38947
rect 2179 38913 2188 38947
rect 2136 38904 2188 38913
rect 1308 38836 1360 38888
rect 1768 38836 1820 38888
rect 5080 38904 5132 38956
rect 10140 38947 10192 38956
rect 10140 38913 10149 38947
rect 10149 38913 10183 38947
rect 10183 38913 10192 38947
rect 10140 38904 10192 38913
rect 3884 38836 3936 38888
rect 9864 38700 9916 38752
rect 2582 38598 2634 38650
rect 2646 38598 2698 38650
rect 2710 38598 2762 38650
rect 2774 38598 2826 38650
rect 2838 38598 2890 38650
rect 5845 38598 5897 38650
rect 5909 38598 5961 38650
rect 5973 38598 6025 38650
rect 6037 38598 6089 38650
rect 6101 38598 6153 38650
rect 9109 38598 9161 38650
rect 9173 38598 9225 38650
rect 9237 38598 9289 38650
rect 9301 38598 9353 38650
rect 9365 38598 9417 38650
rect 2320 38496 2372 38548
rect 3792 38496 3844 38548
rect 7012 38428 7064 38480
rect 1308 38360 1360 38412
rect 1400 38335 1452 38344
rect 1400 38301 1409 38335
rect 1409 38301 1443 38335
rect 1443 38301 1452 38335
rect 1400 38292 1452 38301
rect 2136 38335 2188 38344
rect 2136 38301 2145 38335
rect 2145 38301 2179 38335
rect 2179 38301 2188 38335
rect 2136 38292 2188 38301
rect 2780 38335 2832 38344
rect 2780 38301 2789 38335
rect 2789 38301 2823 38335
rect 2823 38301 2832 38335
rect 2780 38292 2832 38301
rect 756 38156 808 38208
rect 3608 38156 3660 38208
rect 9956 38292 10008 38344
rect 10140 38335 10192 38344
rect 10140 38301 10149 38335
rect 10149 38301 10183 38335
rect 10183 38301 10192 38335
rect 10140 38292 10192 38301
rect 5632 38156 5684 38208
rect 9956 38199 10008 38208
rect 9956 38165 9965 38199
rect 9965 38165 9999 38199
rect 9999 38165 10008 38199
rect 9956 38156 10008 38165
rect 4213 38054 4265 38106
rect 4277 38054 4329 38106
rect 4341 38054 4393 38106
rect 4405 38054 4457 38106
rect 4469 38054 4521 38106
rect 7477 38054 7529 38106
rect 7541 38054 7593 38106
rect 7605 38054 7657 38106
rect 7669 38054 7721 38106
rect 7733 38054 7785 38106
rect 6184 37952 6236 38004
rect 1400 37859 1452 37868
rect 1400 37825 1409 37859
rect 1409 37825 1443 37859
rect 1443 37825 1452 37859
rect 1400 37816 1452 37825
rect 2780 37816 2832 37868
rect 9864 37816 9916 37868
rect 2320 37748 2372 37800
rect 3056 37748 3108 37800
rect 3884 37612 3936 37664
rect 6184 37612 6236 37664
rect 2582 37510 2634 37562
rect 2646 37510 2698 37562
rect 2710 37510 2762 37562
rect 2774 37510 2826 37562
rect 2838 37510 2890 37562
rect 5845 37510 5897 37562
rect 5909 37510 5961 37562
rect 5973 37510 6025 37562
rect 6037 37510 6089 37562
rect 6101 37510 6153 37562
rect 9109 37510 9161 37562
rect 9173 37510 9225 37562
rect 9237 37510 9289 37562
rect 9301 37510 9353 37562
rect 9365 37510 9417 37562
rect 388 37340 440 37392
rect 1308 37340 1360 37392
rect 2320 37272 2372 37324
rect 1400 37247 1452 37256
rect 1400 37213 1409 37247
rect 1409 37213 1443 37247
rect 1443 37213 1452 37247
rect 1400 37204 1452 37213
rect 2688 37247 2740 37256
rect 2688 37213 2697 37247
rect 2697 37213 2731 37247
rect 2731 37213 2740 37247
rect 2688 37204 2740 37213
rect 9956 37204 10008 37256
rect 10140 37247 10192 37256
rect 10140 37213 10149 37247
rect 10149 37213 10183 37247
rect 10183 37213 10192 37247
rect 10140 37204 10192 37213
rect 3056 37136 3108 37188
rect 4988 37136 5040 37188
rect 6460 37068 6512 37120
rect 9956 37111 10008 37120
rect 9956 37077 9965 37111
rect 9965 37077 9999 37111
rect 9999 37077 10008 37111
rect 9956 37068 10008 37077
rect 4213 36966 4265 37018
rect 4277 36966 4329 37018
rect 4341 36966 4393 37018
rect 4405 36966 4457 37018
rect 4469 36966 4521 37018
rect 7477 36966 7529 37018
rect 7541 36966 7593 37018
rect 7605 36966 7657 37018
rect 7669 36966 7721 37018
rect 7733 36966 7785 37018
rect 1952 36864 2004 36916
rect 3700 36864 3752 36916
rect 2688 36796 2740 36848
rect 1400 36771 1452 36780
rect 1400 36737 1409 36771
rect 1409 36737 1443 36771
rect 1443 36737 1452 36771
rect 1400 36728 1452 36737
rect 2136 36771 2188 36780
rect 2136 36737 2145 36771
rect 2145 36737 2179 36771
rect 2179 36737 2188 36771
rect 2136 36728 2188 36737
rect 1124 36660 1176 36712
rect 3792 36796 3844 36848
rect 9956 36728 10008 36780
rect 10140 36771 10192 36780
rect 10140 36737 10149 36771
rect 10149 36737 10183 36771
rect 10183 36737 10192 36771
rect 10140 36728 10192 36737
rect 20 36524 72 36576
rect 756 36524 808 36576
rect 4804 36592 4856 36644
rect 3332 36524 3384 36576
rect 3516 36524 3568 36576
rect 3884 36524 3936 36576
rect 4068 36524 4120 36576
rect 4344 36524 4396 36576
rect 2582 36422 2634 36474
rect 2646 36422 2698 36474
rect 2710 36422 2762 36474
rect 2774 36422 2826 36474
rect 2838 36422 2890 36474
rect 5845 36422 5897 36474
rect 5909 36422 5961 36474
rect 5973 36422 6025 36474
rect 6037 36422 6089 36474
rect 6101 36422 6153 36474
rect 9109 36422 9161 36474
rect 9173 36422 9225 36474
rect 9237 36422 9289 36474
rect 9301 36422 9353 36474
rect 9365 36422 9417 36474
rect 480 36320 532 36372
rect 3608 36320 3660 36372
rect 1492 36252 1544 36304
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 2136 36159 2188 36168
rect 2136 36125 2145 36159
rect 2145 36125 2179 36159
rect 2179 36125 2188 36159
rect 2136 36116 2188 36125
rect 4988 36184 5040 36236
rect 3792 36116 3844 36168
rect 4344 36159 4396 36168
rect 4344 36125 4353 36159
rect 4353 36125 4387 36159
rect 4387 36125 4396 36159
rect 4344 36116 4396 36125
rect 10140 36159 10192 36168
rect 10140 36125 10149 36159
rect 10149 36125 10183 36159
rect 10183 36125 10192 36159
rect 10140 36116 10192 36125
rect 4804 36048 4856 36100
rect 1584 35980 1636 36032
rect 5172 35980 5224 36032
rect 9956 36023 10008 36032
rect 9956 35989 9965 36023
rect 9965 35989 9999 36023
rect 9999 35989 10008 36023
rect 9956 35980 10008 35989
rect 4213 35878 4265 35930
rect 4277 35878 4329 35930
rect 4341 35878 4393 35930
rect 4405 35878 4457 35930
rect 4469 35878 4521 35930
rect 7477 35878 7529 35930
rect 7541 35878 7593 35930
rect 7605 35878 7657 35930
rect 7669 35878 7721 35930
rect 7733 35878 7785 35930
rect 1676 35776 1728 35828
rect 5264 35776 5316 35828
rect 4252 35708 4304 35760
rect 1400 35683 1452 35692
rect 1400 35649 1409 35683
rect 1409 35649 1443 35683
rect 1443 35649 1452 35683
rect 1400 35640 1452 35649
rect 2136 35683 2188 35692
rect 2136 35649 2145 35683
rect 2145 35649 2179 35683
rect 2179 35649 2188 35683
rect 2136 35640 2188 35649
rect 480 35572 532 35624
rect 9956 35640 10008 35692
rect 4620 35572 4672 35624
rect 5448 35572 5500 35624
rect 5540 35504 5592 35556
rect 5172 35436 5224 35488
rect 5356 35436 5408 35488
rect 2582 35334 2634 35386
rect 2646 35334 2698 35386
rect 2710 35334 2762 35386
rect 2774 35334 2826 35386
rect 2838 35334 2890 35386
rect 5845 35334 5897 35386
rect 5909 35334 5961 35386
rect 5973 35334 6025 35386
rect 6037 35334 6089 35386
rect 6101 35334 6153 35386
rect 9109 35334 9161 35386
rect 9173 35334 9225 35386
rect 9237 35334 9289 35386
rect 9301 35334 9353 35386
rect 9365 35334 9417 35386
rect 1216 35232 1268 35284
rect 204 35164 256 35216
rect 3976 35164 4028 35216
rect 1400 35071 1452 35080
rect 1400 35037 1409 35071
rect 1409 35037 1443 35071
rect 1443 35037 1452 35071
rect 1400 35028 1452 35037
rect 10140 35071 10192 35080
rect 1768 34960 1820 35012
rect 4252 34960 4304 35012
rect 4804 34892 4856 34944
rect 10140 35037 10149 35071
rect 10149 35037 10183 35071
rect 10183 35037 10192 35071
rect 10140 35028 10192 35037
rect 4213 34790 4265 34842
rect 4277 34790 4329 34842
rect 4341 34790 4393 34842
rect 4405 34790 4457 34842
rect 4469 34790 4521 34842
rect 7477 34790 7529 34842
rect 7541 34790 7593 34842
rect 7605 34790 7657 34842
rect 7669 34790 7721 34842
rect 7733 34790 7785 34842
rect 4988 34688 5040 34740
rect 5356 34688 5408 34740
rect 6644 34620 6696 34672
rect 1400 34595 1452 34604
rect 1400 34561 1409 34595
rect 1409 34561 1443 34595
rect 1443 34561 1452 34595
rect 1400 34552 1452 34561
rect 3792 34484 3844 34536
rect 4988 34484 5040 34536
rect 10140 34416 10192 34468
rect 2582 34246 2634 34298
rect 2646 34246 2698 34298
rect 2710 34246 2762 34298
rect 2774 34246 2826 34298
rect 2838 34246 2890 34298
rect 5845 34246 5897 34298
rect 5909 34246 5961 34298
rect 5973 34246 6025 34298
rect 6037 34246 6089 34298
rect 6101 34246 6153 34298
rect 9109 34246 9161 34298
rect 9173 34246 9225 34298
rect 9237 34246 9289 34298
rect 9301 34246 9353 34298
rect 9365 34246 9417 34298
rect 5724 34144 5776 34196
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 10140 33983 10192 33992
rect 10140 33949 10149 33983
rect 10149 33949 10183 33983
rect 10183 33949 10192 33983
rect 10140 33940 10192 33949
rect 9864 33804 9916 33856
rect 4213 33702 4265 33754
rect 4277 33702 4329 33754
rect 4341 33702 4393 33754
rect 4405 33702 4457 33754
rect 4469 33702 4521 33754
rect 7477 33702 7529 33754
rect 7541 33702 7593 33754
rect 7605 33702 7657 33754
rect 7669 33702 7721 33754
rect 7733 33702 7785 33754
rect 1584 33643 1636 33652
rect 1584 33609 1593 33643
rect 1593 33609 1627 33643
rect 1627 33609 1636 33643
rect 1584 33600 1636 33609
rect 1400 33507 1452 33516
rect 1400 33473 1409 33507
rect 1409 33473 1443 33507
rect 1443 33473 1452 33507
rect 1400 33464 1452 33473
rect 2582 33158 2634 33210
rect 2646 33158 2698 33210
rect 2710 33158 2762 33210
rect 2774 33158 2826 33210
rect 2838 33158 2890 33210
rect 5845 33158 5897 33210
rect 5909 33158 5961 33210
rect 5973 33158 6025 33210
rect 6037 33158 6089 33210
rect 6101 33158 6153 33210
rect 9109 33158 9161 33210
rect 9173 33158 9225 33210
rect 9237 33158 9289 33210
rect 9301 33158 9353 33210
rect 9365 33158 9417 33210
rect 940 33056 992 33108
rect 1400 32895 1452 32904
rect 1400 32861 1409 32895
rect 1409 32861 1443 32895
rect 1443 32861 1452 32895
rect 1400 32852 1452 32861
rect 10140 32895 10192 32904
rect 10140 32861 10149 32895
rect 10149 32861 10183 32895
rect 10183 32861 10192 32895
rect 10140 32852 10192 32861
rect 9956 32759 10008 32768
rect 9956 32725 9965 32759
rect 9965 32725 9999 32759
rect 9999 32725 10008 32759
rect 9956 32716 10008 32725
rect 4213 32614 4265 32666
rect 4277 32614 4329 32666
rect 4341 32614 4393 32666
rect 4405 32614 4457 32666
rect 4469 32614 4521 32666
rect 7477 32614 7529 32666
rect 7541 32614 7593 32666
rect 7605 32614 7657 32666
rect 7669 32614 7721 32666
rect 7733 32614 7785 32666
rect 1032 32512 1084 32564
rect 2228 32555 2280 32564
rect 2228 32521 2237 32555
rect 2237 32521 2271 32555
rect 2271 32521 2280 32555
rect 2228 32512 2280 32521
rect 1308 32376 1360 32428
rect 2136 32419 2188 32428
rect 2136 32385 2145 32419
rect 2145 32385 2179 32419
rect 2179 32385 2188 32419
rect 2136 32376 2188 32385
rect 3148 32376 3200 32428
rect 10140 32419 10192 32428
rect 10140 32385 10149 32419
rect 10149 32385 10183 32419
rect 10183 32385 10192 32419
rect 10140 32376 10192 32385
rect 1676 32240 1728 32292
rect 6460 32240 6512 32292
rect 9772 32172 9824 32224
rect 2582 32070 2634 32122
rect 2646 32070 2698 32122
rect 2710 32070 2762 32122
rect 2774 32070 2826 32122
rect 2838 32070 2890 32122
rect 5845 32070 5897 32122
rect 5909 32070 5961 32122
rect 5973 32070 6025 32122
rect 6037 32070 6089 32122
rect 6101 32070 6153 32122
rect 9109 32070 9161 32122
rect 9173 32070 9225 32122
rect 9237 32070 9289 32122
rect 9301 32070 9353 32122
rect 9365 32070 9417 32122
rect 2412 31968 2464 32020
rect 3148 31900 3200 31952
rect 5540 31900 5592 31952
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 2136 31807 2188 31816
rect 2136 31773 2145 31807
rect 2145 31773 2179 31807
rect 2179 31773 2188 31807
rect 2136 31764 2188 31773
rect 204 31696 256 31748
rect 9864 31764 9916 31816
rect 3148 31696 3200 31748
rect 4213 31526 4265 31578
rect 4277 31526 4329 31578
rect 4341 31526 4393 31578
rect 4405 31526 4457 31578
rect 4469 31526 4521 31578
rect 7477 31526 7529 31578
rect 7541 31526 7593 31578
rect 7605 31526 7657 31578
rect 7669 31526 7721 31578
rect 7733 31526 7785 31578
rect 1676 31424 1728 31476
rect 2044 31424 2096 31476
rect 3148 31467 3200 31476
rect 3148 31433 3157 31467
rect 3157 31433 3191 31467
rect 3191 31433 3200 31467
rect 3148 31424 3200 31433
rect 1308 31288 1360 31340
rect 2136 31331 2188 31340
rect 2136 31297 2145 31331
rect 2145 31297 2179 31331
rect 2179 31297 2188 31331
rect 2136 31288 2188 31297
rect 3148 31288 3200 31340
rect 9956 31288 10008 31340
rect 10140 31331 10192 31340
rect 10140 31297 10149 31331
rect 10149 31297 10183 31331
rect 10183 31297 10192 31331
rect 10140 31288 10192 31297
rect 1676 31152 1728 31204
rect 8392 31152 8444 31204
rect 3332 31084 3384 31136
rect 4712 31084 4764 31136
rect 9864 31084 9916 31136
rect 2582 30982 2634 31034
rect 2646 30982 2698 31034
rect 2710 30982 2762 31034
rect 2774 30982 2826 31034
rect 2838 30982 2890 31034
rect 5845 30982 5897 31034
rect 5909 30982 5961 31034
rect 5973 30982 6025 31034
rect 6037 30982 6089 31034
rect 6101 30982 6153 31034
rect 9109 30982 9161 31034
rect 9173 30982 9225 31034
rect 9237 30982 9289 31034
rect 9301 30982 9353 31034
rect 9365 30982 9417 31034
rect 1768 30880 1820 30932
rect 2412 30880 2464 30932
rect 2964 30880 3016 30932
rect 4712 30880 4764 30932
rect 5448 30880 5500 30932
rect 940 30812 992 30864
rect 1492 30744 1544 30796
rect 1952 30744 2004 30796
rect 1400 30719 1452 30728
rect 1400 30685 1409 30719
rect 1409 30685 1443 30719
rect 1443 30685 1452 30719
rect 1400 30676 1452 30685
rect 2136 30719 2188 30728
rect 2136 30685 2145 30719
rect 2145 30685 2179 30719
rect 2179 30685 2188 30719
rect 2136 30676 2188 30685
rect 2504 30676 2556 30728
rect 9772 30676 9824 30728
rect 10140 30719 10192 30728
rect 10140 30685 10149 30719
rect 10149 30685 10183 30719
rect 10183 30685 10192 30719
rect 10140 30676 10192 30685
rect 5448 30540 5500 30592
rect 9956 30583 10008 30592
rect 9956 30549 9965 30583
rect 9965 30549 9999 30583
rect 9999 30549 10008 30583
rect 9956 30540 10008 30549
rect 4213 30438 4265 30490
rect 4277 30438 4329 30490
rect 4341 30438 4393 30490
rect 4405 30438 4457 30490
rect 4469 30438 4521 30490
rect 7477 30438 7529 30490
rect 7541 30438 7593 30490
rect 7605 30438 7657 30490
rect 7669 30438 7721 30490
rect 7733 30438 7785 30490
rect 1584 30336 1636 30388
rect 7196 30336 7248 30388
rect 1308 30200 1360 30252
rect 2320 30200 2372 30252
rect 5172 30268 5224 30320
rect 9864 30200 9916 30252
rect 10140 30243 10192 30252
rect 10140 30209 10149 30243
rect 10149 30209 10183 30243
rect 10183 30209 10192 30243
rect 10140 30200 10192 30209
rect 2964 30132 3016 30184
rect 1676 30064 1728 30116
rect 3148 29996 3200 30048
rect 5172 29996 5224 30048
rect 9864 29996 9916 30048
rect 2582 29894 2634 29946
rect 2646 29894 2698 29946
rect 2710 29894 2762 29946
rect 2774 29894 2826 29946
rect 2838 29894 2890 29946
rect 5845 29894 5897 29946
rect 5909 29894 5961 29946
rect 5973 29894 6025 29946
rect 6037 29894 6089 29946
rect 6101 29894 6153 29946
rect 9109 29894 9161 29946
rect 9173 29894 9225 29946
rect 9237 29894 9289 29946
rect 9301 29894 9353 29946
rect 9365 29894 9417 29946
rect 1584 29835 1636 29844
rect 1584 29801 1593 29835
rect 1593 29801 1627 29835
rect 1627 29801 1636 29835
rect 1584 29792 1636 29801
rect 1768 29792 1820 29844
rect 8484 29792 8536 29844
rect 2320 29699 2372 29708
rect 2320 29665 2329 29699
rect 2329 29665 2363 29699
rect 2363 29665 2372 29699
rect 2320 29656 2372 29665
rect 2504 29656 2556 29708
rect 1400 29631 1452 29640
rect 1400 29597 1409 29631
rect 1409 29597 1443 29631
rect 1443 29597 1452 29631
rect 1400 29588 1452 29597
rect 10140 29631 10192 29640
rect 10140 29597 10149 29631
rect 10149 29597 10183 29631
rect 10183 29597 10192 29631
rect 10140 29588 10192 29597
rect 1676 29452 1728 29504
rect 8300 29452 8352 29504
rect 9680 29452 9732 29504
rect 4213 29350 4265 29402
rect 4277 29350 4329 29402
rect 4341 29350 4393 29402
rect 4405 29350 4457 29402
rect 4469 29350 4521 29402
rect 7477 29350 7529 29402
rect 7541 29350 7593 29402
rect 7605 29350 7657 29402
rect 7669 29350 7721 29402
rect 7733 29350 7785 29402
rect 1676 29248 1728 29300
rect 1860 29248 1912 29300
rect 1308 29112 1360 29164
rect 2964 29180 3016 29232
rect 9680 29180 9732 29232
rect 9956 29155 10008 29164
rect 1216 29044 1268 29096
rect 3424 29044 3476 29096
rect 9956 29121 9965 29155
rect 9965 29121 9999 29155
rect 9999 29121 10008 29155
rect 9956 29112 10008 29121
rect 848 28908 900 28960
rect 1492 28908 1544 28960
rect 2044 28908 2096 28960
rect 9956 28976 10008 29028
rect 3424 28908 3476 28960
rect 4712 28908 4764 28960
rect 9864 28951 9916 28960
rect 9864 28917 9873 28951
rect 9873 28917 9907 28951
rect 9907 28917 9916 28951
rect 9864 28908 9916 28917
rect 2582 28806 2634 28858
rect 2646 28806 2698 28858
rect 2710 28806 2762 28858
rect 2774 28806 2826 28858
rect 2838 28806 2890 28858
rect 5845 28806 5897 28858
rect 5909 28806 5961 28858
rect 5973 28806 6025 28858
rect 6037 28806 6089 28858
rect 6101 28806 6153 28858
rect 9109 28806 9161 28858
rect 9173 28806 9225 28858
rect 9237 28806 9289 28858
rect 9301 28806 9353 28858
rect 9365 28806 9417 28858
rect 1952 28704 2004 28756
rect 3884 28704 3936 28756
rect 9956 28747 10008 28756
rect 9956 28713 9965 28747
rect 9965 28713 9999 28747
rect 9999 28713 10008 28747
rect 9956 28704 10008 28713
rect 7012 28636 7064 28688
rect 1400 28543 1452 28552
rect 1400 28509 1409 28543
rect 1409 28509 1443 28543
rect 1443 28509 1452 28543
rect 1400 28500 1452 28509
rect 1032 28364 1084 28416
rect 2872 28500 2924 28552
rect 4712 28500 4764 28552
rect 10140 28543 10192 28552
rect 10140 28509 10149 28543
rect 10149 28509 10183 28543
rect 10183 28509 10192 28543
rect 10140 28500 10192 28509
rect 2504 28364 2556 28416
rect 8760 28364 8812 28416
rect 4213 28262 4265 28314
rect 4277 28262 4329 28314
rect 4341 28262 4393 28314
rect 4405 28262 4457 28314
rect 4469 28262 4521 28314
rect 7477 28262 7529 28314
rect 7541 28262 7593 28314
rect 7605 28262 7657 28314
rect 7669 28262 7721 28314
rect 7733 28262 7785 28314
rect 1768 28160 1820 28212
rect 3516 28160 3568 28212
rect 3884 28160 3936 28212
rect 5080 28160 5132 28212
rect 940 28092 992 28144
rect 1216 28092 1268 28144
rect 1308 28024 1360 28076
rect 1216 27956 1268 28008
rect 2872 28024 2924 28076
rect 10140 28067 10192 28076
rect 10140 28033 10149 28067
rect 10149 28033 10183 28067
rect 10183 28033 10192 28067
rect 10140 28024 10192 28033
rect 4620 27956 4672 28008
rect 1584 27888 1636 27940
rect 9772 27820 9824 27872
rect 2582 27718 2634 27770
rect 2646 27718 2698 27770
rect 2710 27718 2762 27770
rect 2774 27718 2826 27770
rect 2838 27718 2890 27770
rect 5845 27718 5897 27770
rect 5909 27718 5961 27770
rect 5973 27718 6025 27770
rect 6037 27718 6089 27770
rect 6101 27718 6153 27770
rect 9109 27718 9161 27770
rect 9173 27718 9225 27770
rect 9237 27718 9289 27770
rect 9301 27718 9353 27770
rect 9365 27718 9417 27770
rect 2504 27616 2556 27668
rect 2044 27548 2096 27600
rect 3240 27548 3292 27600
rect 3424 27548 3476 27600
rect 4528 27548 4580 27600
rect 664 27480 716 27532
rect 2504 27480 2556 27532
rect 112 27412 164 27464
rect 2320 27412 2372 27464
rect 10232 27412 10284 27464
rect 1952 27387 2004 27396
rect 1952 27353 1961 27387
rect 1961 27353 1995 27387
rect 1995 27353 2004 27387
rect 1952 27344 2004 27353
rect 9864 27276 9916 27328
rect 4213 27174 4265 27226
rect 4277 27174 4329 27226
rect 4341 27174 4393 27226
rect 4405 27174 4457 27226
rect 4469 27174 4521 27226
rect 7477 27174 7529 27226
rect 7541 27174 7593 27226
rect 7605 27174 7657 27226
rect 7669 27174 7721 27226
rect 7733 27174 7785 27226
rect 940 27004 992 27056
rect 1216 27004 1268 27056
rect 10048 26936 10100 26988
rect 9956 26775 10008 26784
rect 9956 26741 9965 26775
rect 9965 26741 9999 26775
rect 9999 26741 10008 26775
rect 9956 26732 10008 26741
rect 2582 26630 2634 26682
rect 2646 26630 2698 26682
rect 2710 26630 2762 26682
rect 2774 26630 2826 26682
rect 2838 26630 2890 26682
rect 5845 26630 5897 26682
rect 5909 26630 5961 26682
rect 5973 26630 6025 26682
rect 6037 26630 6089 26682
rect 6101 26630 6153 26682
rect 9109 26630 9161 26682
rect 9173 26630 9225 26682
rect 9237 26630 9289 26682
rect 9301 26630 9353 26682
rect 9365 26630 9417 26682
rect 8668 26528 8720 26580
rect 9864 26571 9916 26580
rect 9864 26537 9873 26571
rect 9873 26537 9907 26571
rect 9907 26537 9916 26571
rect 9864 26528 9916 26537
rect 10140 26392 10192 26444
rect 9864 26367 9916 26376
rect 9864 26333 9873 26367
rect 9873 26333 9907 26367
rect 9907 26333 9916 26367
rect 9864 26324 9916 26333
rect 1952 26299 2004 26308
rect 1952 26265 1961 26299
rect 1961 26265 1995 26299
rect 1995 26265 2004 26299
rect 1952 26256 2004 26265
rect 4213 26086 4265 26138
rect 4277 26086 4329 26138
rect 4341 26086 4393 26138
rect 4405 26086 4457 26138
rect 4469 26086 4521 26138
rect 7477 26086 7529 26138
rect 7541 26086 7593 26138
rect 7605 26086 7657 26138
rect 7669 26086 7721 26138
rect 7733 26086 7785 26138
rect 8576 25984 8628 26036
rect 10140 26027 10192 26036
rect 10140 25993 10149 26027
rect 10149 25993 10183 26027
rect 10183 25993 10192 26027
rect 10140 25984 10192 25993
rect 9772 25959 9824 25968
rect 9772 25925 9781 25959
rect 9781 25925 9815 25959
rect 9815 25925 9824 25959
rect 9772 25916 9824 25925
rect 9956 25959 10008 25968
rect 9956 25925 9965 25959
rect 9965 25925 9999 25959
rect 9999 25925 10008 25959
rect 9956 25916 10008 25925
rect 1952 25891 2004 25900
rect 1952 25857 1961 25891
rect 1961 25857 1995 25891
rect 1995 25857 2004 25891
rect 1952 25848 2004 25857
rect 2582 25542 2634 25594
rect 2646 25542 2698 25594
rect 2710 25542 2762 25594
rect 2774 25542 2826 25594
rect 2838 25542 2890 25594
rect 5845 25542 5897 25594
rect 5909 25542 5961 25594
rect 5973 25542 6025 25594
rect 6037 25542 6089 25594
rect 6101 25542 6153 25594
rect 9109 25542 9161 25594
rect 9173 25542 9225 25594
rect 9237 25542 9289 25594
rect 9301 25542 9353 25594
rect 9365 25542 9417 25594
rect 7288 25440 7340 25492
rect 10140 25279 10192 25288
rect 10140 25245 10149 25279
rect 10149 25245 10183 25279
rect 10183 25245 10192 25279
rect 10140 25236 10192 25245
rect 1952 25211 2004 25220
rect 1952 25177 1961 25211
rect 1961 25177 1995 25211
rect 1995 25177 2004 25211
rect 1952 25168 2004 25177
rect 9772 25100 9824 25152
rect 4213 24998 4265 25050
rect 4277 24998 4329 25050
rect 4341 24998 4393 25050
rect 4405 24998 4457 25050
rect 4469 24998 4521 25050
rect 7477 24998 7529 25050
rect 7541 24998 7593 25050
rect 7605 24998 7657 25050
rect 7669 24998 7721 25050
rect 7733 24998 7785 25050
rect 1952 24803 2004 24812
rect 1952 24769 1961 24803
rect 1961 24769 1995 24803
rect 1995 24769 2004 24803
rect 1952 24760 2004 24769
rect 2596 24760 2648 24812
rect 3332 24803 3384 24812
rect 2964 24692 3016 24744
rect 3332 24769 3341 24803
rect 3341 24769 3375 24803
rect 3375 24769 3384 24803
rect 3332 24760 3384 24769
rect 10140 24803 10192 24812
rect 10140 24769 10149 24803
rect 10149 24769 10183 24803
rect 10183 24769 10192 24803
rect 10140 24760 10192 24769
rect 7104 24624 7156 24676
rect 2504 24599 2556 24608
rect 2504 24565 2513 24599
rect 2513 24565 2547 24599
rect 2547 24565 2556 24599
rect 2504 24556 2556 24565
rect 3700 24556 3752 24608
rect 9956 24599 10008 24608
rect 9956 24565 9965 24599
rect 9965 24565 9999 24599
rect 9999 24565 10008 24599
rect 9956 24556 10008 24565
rect 2582 24454 2634 24506
rect 2646 24454 2698 24506
rect 2710 24454 2762 24506
rect 2774 24454 2826 24506
rect 2838 24454 2890 24506
rect 5845 24454 5897 24506
rect 5909 24454 5961 24506
rect 5973 24454 6025 24506
rect 6037 24454 6089 24506
rect 6101 24454 6153 24506
rect 9109 24454 9161 24506
rect 9173 24454 9225 24506
rect 9237 24454 9289 24506
rect 9301 24454 9353 24506
rect 9365 24454 9417 24506
rect 1860 24395 1912 24404
rect 1860 24361 1869 24395
rect 1869 24361 1903 24395
rect 1903 24361 1912 24395
rect 1860 24352 1912 24361
rect 1952 24123 2004 24132
rect 1952 24089 1961 24123
rect 1961 24089 1995 24123
rect 1995 24089 2004 24123
rect 1952 24080 2004 24089
rect 6276 24148 6328 24200
rect 10140 24191 10192 24200
rect 10140 24157 10149 24191
rect 10149 24157 10183 24191
rect 10183 24157 10192 24191
rect 10140 24148 10192 24157
rect 2872 24080 2924 24132
rect 1768 24012 1820 24064
rect 9864 24012 9916 24064
rect 4213 23910 4265 23962
rect 4277 23910 4329 23962
rect 4341 23910 4393 23962
rect 4405 23910 4457 23962
rect 4469 23910 4521 23962
rect 7477 23910 7529 23962
rect 7541 23910 7593 23962
rect 7605 23910 7657 23962
rect 7669 23910 7721 23962
rect 7733 23910 7785 23962
rect 2044 23783 2096 23792
rect 2044 23749 2053 23783
rect 2053 23749 2087 23783
rect 2087 23749 2096 23783
rect 2044 23740 2096 23749
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 2872 23672 2924 23724
rect 3056 23672 3108 23724
rect 3608 23715 3660 23724
rect 3608 23681 3617 23715
rect 3617 23681 3651 23715
rect 3651 23681 3660 23715
rect 3608 23672 3660 23681
rect 9956 23715 10008 23724
rect 9956 23681 9965 23715
rect 9965 23681 9999 23715
rect 9999 23681 10008 23715
rect 9956 23672 10008 23681
rect 3792 23604 3844 23656
rect 3332 23536 3384 23588
rect 3148 23468 3200 23520
rect 10140 23468 10192 23520
rect 2582 23366 2634 23418
rect 2646 23366 2698 23418
rect 2710 23366 2762 23418
rect 2774 23366 2826 23418
rect 2838 23366 2890 23418
rect 5845 23366 5897 23418
rect 5909 23366 5961 23418
rect 5973 23366 6025 23418
rect 6037 23366 6089 23418
rect 6101 23366 6153 23418
rect 9109 23366 9161 23418
rect 9173 23366 9225 23418
rect 9237 23366 9289 23418
rect 9301 23366 9353 23418
rect 9365 23366 9417 23418
rect 7840 23264 7892 23316
rect 9864 23307 9916 23316
rect 9864 23273 9873 23307
rect 9873 23273 9907 23307
rect 9907 23273 9916 23307
rect 9864 23264 9916 23273
rect 4896 23128 4948 23180
rect 9772 23171 9824 23180
rect 9772 23137 9781 23171
rect 9781 23137 9815 23171
rect 9815 23137 9824 23171
rect 9772 23128 9824 23137
rect 10048 23128 10100 23180
rect 3792 23103 3844 23112
rect 1952 23035 2004 23044
rect 1952 23001 1961 23035
rect 1961 23001 1995 23035
rect 1995 23001 2004 23035
rect 1952 22992 2004 23001
rect 3792 23069 3801 23103
rect 3801 23069 3835 23103
rect 3835 23069 3844 23103
rect 3792 23060 3844 23069
rect 3976 23103 4028 23112
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 9128 23103 9180 23112
rect 9128 23069 9137 23103
rect 9137 23069 9171 23103
rect 9171 23069 9180 23103
rect 9128 23060 9180 23069
rect 2964 22992 3016 23044
rect 1676 22924 1728 22976
rect 3056 22924 3108 22976
rect 9588 22924 9640 22976
rect 9864 22924 9916 22976
rect 9956 22924 10008 22976
rect 4213 22822 4265 22874
rect 4277 22822 4329 22874
rect 4341 22822 4393 22874
rect 4405 22822 4457 22874
rect 4469 22822 4521 22874
rect 7477 22822 7529 22874
rect 7541 22822 7593 22874
rect 7605 22822 7657 22874
rect 7669 22822 7721 22874
rect 7733 22822 7785 22874
rect 7380 22720 7432 22772
rect 9680 22763 9732 22772
rect 9680 22729 9689 22763
rect 9689 22729 9723 22763
rect 9723 22729 9732 22763
rect 9680 22720 9732 22729
rect 1952 22627 2004 22636
rect 1952 22593 1961 22627
rect 1961 22593 1995 22627
rect 1995 22593 2004 22627
rect 1952 22584 2004 22593
rect 3240 22584 3292 22636
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 9956 22627 10008 22636
rect 9956 22593 9965 22627
rect 9965 22593 9999 22627
rect 9999 22593 10008 22627
rect 9956 22584 10008 22593
rect 10140 22627 10192 22636
rect 10140 22593 10149 22627
rect 10149 22593 10183 22627
rect 10183 22593 10192 22627
rect 10140 22584 10192 22593
rect 2964 22559 3016 22568
rect 2964 22525 2973 22559
rect 2973 22525 3007 22559
rect 3007 22525 3016 22559
rect 2964 22516 3016 22525
rect 9036 22423 9088 22432
rect 9036 22389 9045 22423
rect 9045 22389 9079 22423
rect 9079 22389 9088 22423
rect 9036 22380 9088 22389
rect 2582 22278 2634 22330
rect 2646 22278 2698 22330
rect 2710 22278 2762 22330
rect 2774 22278 2826 22330
rect 2838 22278 2890 22330
rect 5845 22278 5897 22330
rect 5909 22278 5961 22330
rect 5973 22278 6025 22330
rect 6037 22278 6089 22330
rect 6101 22278 6153 22330
rect 9109 22278 9161 22330
rect 9173 22278 9225 22330
rect 9237 22278 9289 22330
rect 9301 22278 9353 22330
rect 9365 22278 9417 22330
rect 8024 22040 8076 22092
rect 9496 22083 9548 22092
rect 9496 22049 9505 22083
rect 9505 22049 9539 22083
rect 9539 22049 9548 22083
rect 9496 22040 9548 22049
rect 1952 22015 2004 22024
rect 1952 21981 1961 22015
rect 1961 21981 1995 22015
rect 1995 21981 2004 22015
rect 1952 21972 2004 21981
rect 2688 22015 2740 22024
rect 2688 21981 2691 22015
rect 2691 21981 2725 22015
rect 2725 21981 2740 22015
rect 2688 21972 2740 21981
rect 3608 21972 3660 22024
rect 9680 21972 9732 22024
rect 9864 22015 9916 22024
rect 9864 21981 9873 22015
rect 9873 21981 9907 22015
rect 9907 21981 9916 22015
rect 9864 21972 9916 21981
rect 10048 22015 10100 22024
rect 10048 21981 10057 22015
rect 10057 21981 10091 22015
rect 10091 21981 10100 22015
rect 10048 21972 10100 21981
rect 2964 21904 3016 21956
rect 3792 21904 3844 21956
rect 1952 21836 2004 21888
rect 3976 21836 4028 21888
rect 4213 21734 4265 21786
rect 4277 21734 4329 21786
rect 4341 21734 4393 21786
rect 4405 21734 4457 21786
rect 4469 21734 4521 21786
rect 7477 21734 7529 21786
rect 7541 21734 7593 21786
rect 7605 21734 7657 21786
rect 7669 21734 7721 21786
rect 7733 21734 7785 21786
rect 572 21632 624 21684
rect 3608 21632 3660 21684
rect 10048 21632 10100 21684
rect 1492 21564 1544 21616
rect 2688 21564 2740 21616
rect 3976 21607 4028 21616
rect 3976 21573 3985 21607
rect 3985 21573 4019 21607
rect 4019 21573 4028 21607
rect 3976 21564 4028 21573
rect 3148 21496 3200 21548
rect 8944 21539 8996 21548
rect 8944 21505 8953 21539
rect 8953 21505 8987 21539
rect 8987 21505 8996 21539
rect 8944 21496 8996 21505
rect 9772 21496 9824 21548
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 1492 21403 1544 21412
rect 1492 21369 1501 21403
rect 1501 21369 1535 21403
rect 1535 21369 1544 21403
rect 1492 21360 1544 21369
rect 2964 21292 3016 21344
rect 3148 21335 3200 21344
rect 3148 21301 3157 21335
rect 3157 21301 3191 21335
rect 3191 21301 3200 21335
rect 3148 21292 3200 21301
rect 3240 21292 3292 21344
rect 3608 21292 3660 21344
rect 9588 21292 9640 21344
rect 9864 21335 9916 21344
rect 9864 21301 9873 21335
rect 9873 21301 9907 21335
rect 9907 21301 9916 21335
rect 9864 21292 9916 21301
rect 2582 21190 2634 21242
rect 2646 21190 2698 21242
rect 2710 21190 2762 21242
rect 2774 21190 2826 21242
rect 2838 21190 2890 21242
rect 5845 21190 5897 21242
rect 5909 21190 5961 21242
rect 5973 21190 6025 21242
rect 6037 21190 6089 21242
rect 6101 21190 6153 21242
rect 9109 21190 9161 21242
rect 9173 21190 9225 21242
rect 9237 21190 9289 21242
rect 9301 21190 9353 21242
rect 9365 21190 9417 21242
rect 9956 21088 10008 21140
rect 9588 20952 9640 21004
rect 3056 20884 3108 20936
rect 9036 20927 9088 20936
rect 9036 20893 9045 20927
rect 9045 20893 9079 20927
rect 9079 20893 9088 20927
rect 9036 20884 9088 20893
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 9680 20884 9732 20893
rect 10140 20884 10192 20936
rect 756 20816 808 20868
rect 2412 20816 2464 20868
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 4213 20646 4265 20698
rect 4277 20646 4329 20698
rect 4341 20646 4393 20698
rect 4405 20646 4457 20698
rect 4469 20646 4521 20698
rect 7477 20646 7529 20698
rect 7541 20646 7593 20698
rect 7605 20646 7657 20698
rect 7669 20646 7721 20698
rect 7733 20646 7785 20698
rect 10048 20544 10100 20596
rect 9128 20476 9180 20528
rect 1952 20408 2004 20460
rect 9956 20451 10008 20460
rect 9956 20417 9965 20451
rect 9965 20417 9999 20451
rect 9999 20417 10008 20451
rect 9956 20408 10008 20417
rect 1492 20315 1544 20324
rect 1492 20281 1501 20315
rect 1501 20281 1535 20315
rect 1535 20281 1544 20315
rect 1492 20272 1544 20281
rect 2582 20102 2634 20154
rect 2646 20102 2698 20154
rect 2710 20102 2762 20154
rect 2774 20102 2826 20154
rect 2838 20102 2890 20154
rect 5845 20102 5897 20154
rect 5909 20102 5961 20154
rect 5973 20102 6025 20154
rect 6037 20102 6089 20154
rect 6101 20102 6153 20154
rect 9109 20102 9161 20154
rect 9173 20102 9225 20154
rect 9237 20102 9289 20154
rect 9301 20102 9353 20154
rect 9365 20102 9417 20154
rect 9956 20043 10008 20052
rect 9956 20009 9965 20043
rect 9965 20009 9999 20043
rect 9999 20009 10008 20043
rect 9956 20000 10008 20009
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 10140 19839 10192 19848
rect 10140 19805 10149 19839
rect 10149 19805 10183 19839
rect 10183 19805 10192 19839
rect 10140 19796 10192 19805
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 4213 19558 4265 19610
rect 4277 19558 4329 19610
rect 4341 19558 4393 19610
rect 4405 19558 4457 19610
rect 4469 19558 4521 19610
rect 7477 19558 7529 19610
rect 7541 19558 7593 19610
rect 7605 19558 7657 19610
rect 7669 19558 7721 19610
rect 7733 19558 7785 19610
rect 9864 19456 9916 19508
rect 296 19388 348 19440
rect 2044 19388 2096 19440
rect 3332 19320 3384 19372
rect 10232 19252 10284 19304
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 2582 19014 2634 19066
rect 2646 19014 2698 19066
rect 2710 19014 2762 19066
rect 2774 19014 2826 19066
rect 2838 19014 2890 19066
rect 5845 19014 5897 19066
rect 5909 19014 5961 19066
rect 5973 19014 6025 19066
rect 6037 19014 6089 19066
rect 6101 19014 6153 19066
rect 9109 19014 9161 19066
rect 9173 19014 9225 19066
rect 9237 19014 9289 19066
rect 9301 19014 9353 19066
rect 9365 19014 9417 19066
rect 1768 18708 1820 18760
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 4213 18470 4265 18522
rect 4277 18470 4329 18522
rect 4341 18470 4393 18522
rect 4405 18470 4457 18522
rect 4469 18470 4521 18522
rect 7477 18470 7529 18522
rect 7541 18470 7593 18522
rect 7605 18470 7657 18522
rect 7669 18470 7721 18522
rect 7733 18470 7785 18522
rect 3792 18300 3844 18352
rect 2320 18275 2372 18284
rect 2320 18241 2329 18275
rect 2329 18241 2363 18275
rect 2363 18241 2372 18275
rect 2320 18232 2372 18241
rect 2228 18164 2280 18216
rect 388 18096 440 18148
rect 2320 18096 2372 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 1676 18028 1728 18080
rect 2964 18028 3016 18080
rect 6736 18028 6788 18080
rect 2582 17926 2634 17978
rect 2646 17926 2698 17978
rect 2710 17926 2762 17978
rect 2774 17926 2826 17978
rect 2838 17926 2890 17978
rect 5845 17926 5897 17978
rect 5909 17926 5961 17978
rect 5973 17926 6025 17978
rect 6037 17926 6089 17978
rect 6101 17926 6153 17978
rect 9109 17926 9161 17978
rect 9173 17926 9225 17978
rect 9237 17926 9289 17978
rect 9301 17926 9353 17978
rect 9365 17926 9417 17978
rect 1952 17824 2004 17876
rect 4068 17824 4120 17876
rect 2504 17688 2556 17740
rect 2228 17620 2280 17672
rect 7932 17620 7984 17672
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 1768 17484 1820 17536
rect 4213 17382 4265 17434
rect 4277 17382 4329 17434
rect 4341 17382 4393 17434
rect 4405 17382 4457 17434
rect 4469 17382 4521 17434
rect 7477 17382 7529 17434
rect 7541 17382 7593 17434
rect 7605 17382 7657 17434
rect 7669 17382 7721 17434
rect 7733 17382 7785 17434
rect 3332 17280 3384 17332
rect 5264 17280 5316 17332
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 2228 17144 2280 17196
rect 6368 17144 6420 17196
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 1676 16940 1728 16992
rect 2582 16838 2634 16890
rect 2646 16838 2698 16890
rect 2710 16838 2762 16890
rect 2774 16838 2826 16890
rect 2838 16838 2890 16890
rect 5845 16838 5897 16890
rect 5909 16838 5961 16890
rect 5973 16838 6025 16890
rect 6037 16838 6089 16890
rect 6101 16838 6153 16890
rect 9109 16838 9161 16890
rect 9173 16838 9225 16890
rect 9237 16838 9289 16890
rect 9301 16838 9353 16890
rect 9365 16838 9417 16890
rect 1860 16668 1912 16720
rect 1768 16532 1820 16584
rect 2228 16600 2280 16652
rect 3792 16736 3844 16788
rect 2964 16668 3016 16720
rect 2412 16532 2464 16584
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 2964 16396 3016 16448
rect 4213 16294 4265 16346
rect 4277 16294 4329 16346
rect 4341 16294 4393 16346
rect 4405 16294 4457 16346
rect 4469 16294 4521 16346
rect 7477 16294 7529 16346
rect 7541 16294 7593 16346
rect 7605 16294 7657 16346
rect 7669 16294 7721 16346
rect 7733 16294 7785 16346
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 6552 16124 6604 16176
rect 3700 16056 3752 16108
rect 3240 15988 3292 16040
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 1676 15852 1728 15904
rect 3056 15852 3108 15904
rect 2582 15750 2634 15802
rect 2646 15750 2698 15802
rect 2710 15750 2762 15802
rect 2774 15750 2826 15802
rect 2838 15750 2890 15802
rect 5845 15750 5897 15802
rect 5909 15750 5961 15802
rect 5973 15750 6025 15802
rect 6037 15750 6089 15802
rect 6101 15750 6153 15802
rect 9109 15750 9161 15802
rect 9173 15750 9225 15802
rect 9237 15750 9289 15802
rect 9301 15750 9353 15802
rect 9365 15750 9417 15802
rect 2964 15580 3016 15632
rect 2044 15512 2096 15564
rect 2136 15487 2188 15496
rect 2136 15453 2145 15487
rect 2145 15453 2179 15487
rect 2179 15453 2188 15487
rect 2136 15444 2188 15453
rect 3240 15512 3292 15564
rect 3424 15512 3476 15564
rect 6828 15444 6880 15496
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 2228 15351 2280 15360
rect 2228 15317 2237 15351
rect 2237 15317 2271 15351
rect 2271 15317 2280 15351
rect 2228 15308 2280 15317
rect 3240 15308 3292 15360
rect 4213 15206 4265 15258
rect 4277 15206 4329 15258
rect 4341 15206 4393 15258
rect 4405 15206 4457 15258
rect 4469 15206 4521 15258
rect 7477 15206 7529 15258
rect 7541 15206 7593 15258
rect 7605 15206 7657 15258
rect 7669 15206 7721 15258
rect 7733 15206 7785 15258
rect 1860 14968 1912 15020
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 3516 15036 3568 15088
rect 3332 14968 3384 15020
rect 3424 15011 3476 15020
rect 3424 14977 3433 15011
rect 3433 14977 3467 15011
rect 3467 14977 3476 15011
rect 3424 14968 3476 14977
rect 6184 14900 6236 14952
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 1768 14764 1820 14816
rect 3056 14764 3108 14816
rect 3424 14807 3476 14816
rect 3424 14773 3433 14807
rect 3433 14773 3467 14807
rect 3467 14773 3476 14807
rect 3424 14764 3476 14773
rect 2582 14662 2634 14714
rect 2646 14662 2698 14714
rect 2710 14662 2762 14714
rect 2774 14662 2826 14714
rect 2838 14662 2890 14714
rect 5845 14662 5897 14714
rect 5909 14662 5961 14714
rect 5973 14662 6025 14714
rect 6037 14662 6089 14714
rect 6101 14662 6153 14714
rect 9109 14662 9161 14714
rect 9173 14662 9225 14714
rect 9237 14662 9289 14714
rect 9301 14662 9353 14714
rect 9365 14662 9417 14714
rect 2964 14492 3016 14544
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 2320 14399 2372 14408
rect 2320 14365 2329 14399
rect 2329 14365 2363 14399
rect 2363 14365 2372 14399
rect 2320 14356 2372 14365
rect 2504 14356 2556 14408
rect 5632 14424 5684 14476
rect 3332 14356 3384 14408
rect 3884 14356 3936 14408
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2136 14220 2188 14272
rect 2964 14220 3016 14272
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 3884 14220 3936 14229
rect 4213 14118 4265 14170
rect 4277 14118 4329 14170
rect 4341 14118 4393 14170
rect 4405 14118 4457 14170
rect 4469 14118 4521 14170
rect 7477 14118 7529 14170
rect 7541 14118 7593 14170
rect 7605 14118 7657 14170
rect 7669 14118 7721 14170
rect 7733 14118 7785 14170
rect 3884 13880 3936 13932
rect 3332 13812 3384 13864
rect 3608 13812 3660 13864
rect 480 13744 532 13796
rect 1400 13744 1452 13796
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 2582 13574 2634 13626
rect 2646 13574 2698 13626
rect 2710 13574 2762 13626
rect 2774 13574 2826 13626
rect 2838 13574 2890 13626
rect 5845 13574 5897 13626
rect 5909 13574 5961 13626
rect 5973 13574 6025 13626
rect 6037 13574 6089 13626
rect 6101 13574 6153 13626
rect 9109 13574 9161 13626
rect 9173 13574 9225 13626
rect 9237 13574 9289 13626
rect 9301 13574 9353 13626
rect 9365 13574 9417 13626
rect 2504 13472 2556 13524
rect 3424 13404 3476 13456
rect 2780 13268 2832 13320
rect 3608 13268 3660 13320
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 4213 13030 4265 13082
rect 4277 13030 4329 13082
rect 4341 13030 4393 13082
rect 4405 13030 4457 13082
rect 4469 13030 4521 13082
rect 7477 13030 7529 13082
rect 7541 13030 7593 13082
rect 7605 13030 7657 13082
rect 7669 13030 7721 13082
rect 7733 13030 7785 13082
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 2780 12792 2832 12844
rect 3792 12792 3844 12844
rect 1124 12724 1176 12776
rect 3332 12724 3384 12776
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 3976 12588 4028 12640
rect 5448 12588 5500 12640
rect 2582 12486 2634 12538
rect 2646 12486 2698 12538
rect 2710 12486 2762 12538
rect 2774 12486 2826 12538
rect 2838 12486 2890 12538
rect 5845 12486 5897 12538
rect 5909 12486 5961 12538
rect 5973 12486 6025 12538
rect 6037 12486 6089 12538
rect 6101 12486 6153 12538
rect 9109 12486 9161 12538
rect 9173 12486 9225 12538
rect 9237 12486 9289 12538
rect 9301 12486 9353 12538
rect 9365 12486 9417 12538
rect 204 12384 256 12436
rect 1584 12384 1636 12436
rect 3240 12180 3292 12232
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 4213 11942 4265 11994
rect 4277 11942 4329 11994
rect 4341 11942 4393 11994
rect 4405 11942 4457 11994
rect 4469 11942 4521 11994
rect 7477 11942 7529 11994
rect 7541 11942 7593 11994
rect 7605 11942 7657 11994
rect 7669 11942 7721 11994
rect 7733 11942 7785 11994
rect 3056 11704 3108 11756
rect 1492 11543 1544 11552
rect 1492 11509 1501 11543
rect 1501 11509 1535 11543
rect 1535 11509 1544 11543
rect 1492 11500 1544 11509
rect 2582 11398 2634 11450
rect 2646 11398 2698 11450
rect 2710 11398 2762 11450
rect 2774 11398 2826 11450
rect 2838 11398 2890 11450
rect 5845 11398 5897 11450
rect 5909 11398 5961 11450
rect 5973 11398 6025 11450
rect 6037 11398 6089 11450
rect 6101 11398 6153 11450
rect 9109 11398 9161 11450
rect 9173 11398 9225 11450
rect 9237 11398 9289 11450
rect 9301 11398 9353 11450
rect 9365 11398 9417 11450
rect 2228 11092 2280 11144
rect 3424 11024 3476 11076
rect 5172 11024 5224 11076
rect 1492 10999 1544 11008
rect 1492 10965 1501 10999
rect 1501 10965 1535 10999
rect 1535 10965 1544 10999
rect 1492 10956 1544 10965
rect 4213 10854 4265 10906
rect 4277 10854 4329 10906
rect 4341 10854 4393 10906
rect 4405 10854 4457 10906
rect 4469 10854 4521 10906
rect 7477 10854 7529 10906
rect 7541 10854 7593 10906
rect 7605 10854 7657 10906
rect 7669 10854 7721 10906
rect 7733 10854 7785 10906
rect 2964 10616 3016 10668
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 2582 10310 2634 10362
rect 2646 10310 2698 10362
rect 2710 10310 2762 10362
rect 2774 10310 2826 10362
rect 2838 10310 2890 10362
rect 5845 10310 5897 10362
rect 5909 10310 5961 10362
rect 5973 10310 6025 10362
rect 6037 10310 6089 10362
rect 6101 10310 6153 10362
rect 9109 10310 9161 10362
rect 9173 10310 9225 10362
rect 9237 10310 9289 10362
rect 9301 10310 9353 10362
rect 9365 10310 9417 10362
rect 3608 10072 3660 10124
rect 1768 10004 1820 10056
rect 3056 10004 3108 10056
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 4213 9766 4265 9818
rect 4277 9766 4329 9818
rect 4341 9766 4393 9818
rect 4405 9766 4457 9818
rect 4469 9766 4521 9818
rect 7477 9766 7529 9818
rect 7541 9766 7593 9818
rect 7605 9766 7657 9818
rect 7669 9766 7721 9818
rect 7733 9766 7785 9818
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 1492 9367 1544 9376
rect 1492 9333 1501 9367
rect 1501 9333 1535 9367
rect 1535 9333 1544 9367
rect 1492 9324 1544 9333
rect 2320 9367 2372 9376
rect 2320 9333 2329 9367
rect 2329 9333 2363 9367
rect 2363 9333 2372 9367
rect 2320 9324 2372 9333
rect 2582 9222 2634 9274
rect 2646 9222 2698 9274
rect 2710 9222 2762 9274
rect 2774 9222 2826 9274
rect 2838 9222 2890 9274
rect 5845 9222 5897 9274
rect 5909 9222 5961 9274
rect 5973 9222 6025 9274
rect 6037 9222 6089 9274
rect 6101 9222 6153 9274
rect 9109 9222 9161 9274
rect 9173 9222 9225 9274
rect 9237 9222 9289 9274
rect 9301 9222 9353 9274
rect 9365 9222 9417 9274
rect 1676 9120 1728 9172
rect 940 9052 992 9104
rect 2320 9052 2372 9104
rect 1400 8984 1452 9036
rect 2228 8916 2280 8968
rect 3056 8916 3108 8968
rect 3332 8916 3384 8968
rect 1400 8780 1452 8832
rect 1676 8780 1728 8832
rect 4213 8678 4265 8730
rect 4277 8678 4329 8730
rect 4341 8678 4393 8730
rect 4405 8678 4457 8730
rect 4469 8678 4521 8730
rect 7477 8678 7529 8730
rect 7541 8678 7593 8730
rect 7605 8678 7657 8730
rect 7669 8678 7721 8730
rect 7733 8678 7785 8730
rect 2228 8576 2280 8628
rect 1584 8508 1636 8560
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 3056 8508 3108 8560
rect 3516 8440 3568 8492
rect 4988 8440 5040 8492
rect 5356 8372 5408 8424
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 1676 8304 1728 8356
rect 2964 8236 3016 8288
rect 2582 8134 2634 8186
rect 2646 8134 2698 8186
rect 2710 8134 2762 8186
rect 2774 8134 2826 8186
rect 2838 8134 2890 8186
rect 5845 8134 5897 8186
rect 5909 8134 5961 8186
rect 5973 8134 6025 8186
rect 6037 8134 6089 8186
rect 6101 8134 6153 8186
rect 9109 8134 9161 8186
rect 9173 8134 9225 8186
rect 9237 8134 9289 8186
rect 9301 8134 9353 8186
rect 9365 8134 9417 8186
rect 2964 7964 3016 8016
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 5540 7896 5592 7948
rect 3516 7828 3568 7880
rect 4804 7828 4856 7880
rect 3240 7760 3292 7812
rect 1308 7692 1360 7744
rect 2228 7735 2280 7744
rect 2228 7701 2237 7735
rect 2237 7701 2271 7735
rect 2271 7701 2280 7735
rect 2228 7692 2280 7701
rect 2964 7692 3016 7744
rect 3056 7692 3108 7744
rect 4213 7590 4265 7642
rect 4277 7590 4329 7642
rect 4341 7590 4393 7642
rect 4405 7590 4457 7642
rect 4469 7590 4521 7642
rect 7477 7590 7529 7642
rect 7541 7590 7593 7642
rect 7605 7590 7657 7642
rect 7669 7590 7721 7642
rect 7733 7590 7785 7642
rect 1952 7488 2004 7540
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 3056 7352 3108 7404
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 3424 7395 3476 7404
rect 3424 7361 3433 7395
rect 3433 7361 3467 7395
rect 3467 7361 3476 7395
rect 3424 7352 3476 7361
rect 2044 7148 2096 7200
rect 3332 7148 3384 7200
rect 2582 7046 2634 7098
rect 2646 7046 2698 7098
rect 2710 7046 2762 7098
rect 2774 7046 2826 7098
rect 2838 7046 2890 7098
rect 5845 7046 5897 7098
rect 5909 7046 5961 7098
rect 5973 7046 6025 7098
rect 6037 7046 6089 7098
rect 6101 7046 6153 7098
rect 9109 7046 9161 7098
rect 9173 7046 9225 7098
rect 9237 7046 9289 7098
rect 9301 7046 9353 7098
rect 9365 7046 9417 7098
rect 2964 6808 3016 6860
rect 3148 6851 3200 6860
rect 3148 6817 3157 6851
rect 3157 6817 3191 6851
rect 3191 6817 3200 6851
rect 3148 6808 3200 6817
rect 3976 6783 4028 6792
rect 3240 6672 3292 6724
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 1492 6647 1544 6656
rect 1492 6613 1501 6647
rect 1501 6613 1535 6647
rect 1535 6613 1544 6647
rect 1492 6604 1544 6613
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 9956 6647 10008 6656
rect 9956 6613 9965 6647
rect 9965 6613 9999 6647
rect 9999 6613 10008 6647
rect 9956 6604 10008 6613
rect 4213 6502 4265 6554
rect 4277 6502 4329 6554
rect 4341 6502 4393 6554
rect 4405 6502 4457 6554
rect 4469 6502 4521 6554
rect 7477 6502 7529 6554
rect 7541 6502 7593 6554
rect 7605 6502 7657 6554
rect 7669 6502 7721 6554
rect 7733 6502 7785 6554
rect 2320 6400 2372 6452
rect 9956 6332 10008 6384
rect 3148 6264 3200 6316
rect 2964 6239 3016 6248
rect 2964 6205 2973 6239
rect 2973 6205 3007 6239
rect 3007 6205 3016 6239
rect 2964 6196 3016 6205
rect 9956 6196 10008 6248
rect 1124 6128 1176 6180
rect 2582 5958 2634 6010
rect 2646 5958 2698 6010
rect 2710 5958 2762 6010
rect 2774 5958 2826 6010
rect 2838 5958 2890 6010
rect 5845 5958 5897 6010
rect 5909 5958 5961 6010
rect 5973 5958 6025 6010
rect 6037 5958 6089 6010
rect 6101 5958 6153 6010
rect 9109 5958 9161 6010
rect 9173 5958 9225 6010
rect 9237 5958 9289 6010
rect 9301 5958 9353 6010
rect 9365 5958 9417 6010
rect 4620 5856 4672 5908
rect 4712 5899 4764 5908
rect 4712 5865 4721 5899
rect 4721 5865 4755 5899
rect 4755 5865 4764 5899
rect 4712 5856 4764 5865
rect 1032 5720 1084 5772
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 2044 5652 2096 5704
rect 9864 5652 9916 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2136 5516 2188 5568
rect 4213 5414 4265 5466
rect 4277 5414 4329 5466
rect 4341 5414 4393 5466
rect 4405 5414 4457 5466
rect 4469 5414 4521 5466
rect 7477 5414 7529 5466
rect 7541 5414 7593 5466
rect 7605 5414 7657 5466
rect 7669 5414 7721 5466
rect 7733 5414 7785 5466
rect 3884 5312 3936 5364
rect 9956 5355 10008 5364
rect 9956 5321 9965 5355
rect 9965 5321 9999 5355
rect 9999 5321 10008 5355
rect 9956 5312 10008 5321
rect 2044 5244 2096 5296
rect 2596 5244 2648 5296
rect 2872 5176 2924 5228
rect 3056 5176 3108 5228
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 10140 5219 10192 5228
rect 10140 5185 10149 5219
rect 10149 5185 10183 5219
rect 10183 5185 10192 5219
rect 10140 5176 10192 5185
rect 4712 5108 4764 5160
rect 3148 5040 3200 5092
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 2964 4972 3016 5024
rect 2582 4870 2634 4922
rect 2646 4870 2698 4922
rect 2710 4870 2762 4922
rect 2774 4870 2826 4922
rect 2838 4870 2890 4922
rect 5845 4870 5897 4922
rect 5909 4870 5961 4922
rect 5973 4870 6025 4922
rect 6037 4870 6089 4922
rect 6101 4870 6153 4922
rect 9109 4870 9161 4922
rect 9173 4870 9225 4922
rect 9237 4870 9289 4922
rect 9301 4870 9353 4922
rect 9365 4870 9417 4922
rect 1216 4768 1268 4820
rect 3056 4768 3108 4820
rect 3332 4700 3384 4752
rect 1124 4496 1176 4548
rect 2504 4564 2556 4616
rect 4620 4564 4672 4616
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 1676 4428 1728 4480
rect 2872 4471 2924 4480
rect 2872 4437 2881 4471
rect 2881 4437 2915 4471
rect 2915 4437 2924 4471
rect 2872 4428 2924 4437
rect 4213 4326 4265 4378
rect 4277 4326 4329 4378
rect 4341 4326 4393 4378
rect 4405 4326 4457 4378
rect 4469 4326 4521 4378
rect 7477 4326 7529 4378
rect 7541 4326 7593 4378
rect 7605 4326 7657 4378
rect 7669 4326 7721 4378
rect 7733 4326 7785 4378
rect 4068 4224 4120 4276
rect 2228 4088 2280 4140
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 2872 4020 2924 4072
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 2320 3884 2372 3893
rect 2582 3782 2634 3834
rect 2646 3782 2698 3834
rect 2710 3782 2762 3834
rect 2774 3782 2826 3834
rect 2838 3782 2890 3834
rect 5845 3782 5897 3834
rect 5909 3782 5961 3834
rect 5973 3782 6025 3834
rect 6037 3782 6089 3834
rect 6101 3782 6153 3834
rect 9109 3782 9161 3834
rect 9173 3782 9225 3834
rect 9237 3782 9289 3834
rect 9301 3782 9353 3834
rect 9365 3782 9417 3834
rect 9864 3680 9916 3732
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 1952 3476 2004 3528
rect 9864 3476 9916 3528
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 1400 3340 1452 3392
rect 1676 3340 1728 3392
rect 4213 3238 4265 3290
rect 4277 3238 4329 3290
rect 4341 3238 4393 3290
rect 4405 3238 4457 3290
rect 4469 3238 4521 3290
rect 7477 3238 7529 3290
rect 7541 3238 7593 3290
rect 7605 3238 7657 3290
rect 7669 3238 7721 3290
rect 7733 3238 7785 3290
rect 2964 3000 3016 3052
rect 9864 3043 9916 3052
rect 9864 3009 9873 3043
rect 9873 3009 9907 3043
rect 9907 3009 9916 3043
rect 9864 3000 9916 3009
rect 10140 2975 10192 2984
rect 10140 2941 10149 2975
rect 10149 2941 10183 2975
rect 10183 2941 10192 2975
rect 10140 2932 10192 2941
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 2582 2694 2634 2746
rect 2646 2694 2698 2746
rect 2710 2694 2762 2746
rect 2774 2694 2826 2746
rect 2838 2694 2890 2746
rect 5845 2694 5897 2746
rect 5909 2694 5961 2746
rect 5973 2694 6025 2746
rect 6037 2694 6089 2746
rect 6101 2694 6153 2746
rect 9109 2694 9161 2746
rect 9173 2694 9225 2746
rect 9237 2694 9289 2746
rect 9301 2694 9353 2746
rect 9365 2694 9417 2746
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 2964 2388 3016 2440
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 1400 2252 1452 2304
rect 2780 2252 2832 2304
rect 3056 2295 3108 2304
rect 3056 2261 3065 2295
rect 3065 2261 3099 2295
rect 3099 2261 3108 2295
rect 3056 2252 3108 2261
rect 4213 2150 4265 2202
rect 4277 2150 4329 2202
rect 4341 2150 4393 2202
rect 4405 2150 4457 2202
rect 4469 2150 4521 2202
rect 7477 2150 7529 2202
rect 7541 2150 7593 2202
rect 7605 2150 7657 2202
rect 7669 2150 7721 2202
rect 7733 2150 7785 2202
<< metal2 >>
rect 3790 79656 3846 79665
rect 3790 79591 3846 79600
rect 3054 79112 3110 79121
rect 3054 79047 3110 79056
rect 1490 78568 1546 78577
rect 1490 78503 1546 78512
rect 1400 77512 1452 77518
rect 1400 77454 1452 77460
rect 1308 77036 1360 77042
rect 1308 76978 1360 76984
rect 1320 76401 1348 76978
rect 1412 76945 1440 77454
rect 1504 77042 1532 78503
rect 2962 78024 3018 78033
rect 2962 77959 3018 77968
rect 2582 77820 2890 77840
rect 2582 77818 2588 77820
rect 2644 77818 2668 77820
rect 2724 77818 2748 77820
rect 2804 77818 2828 77820
rect 2884 77818 2890 77820
rect 2644 77766 2646 77818
rect 2826 77766 2828 77818
rect 2582 77764 2588 77766
rect 2644 77764 2668 77766
rect 2724 77764 2748 77766
rect 2804 77764 2828 77766
rect 2884 77764 2890 77766
rect 2582 77744 2890 77764
rect 1768 77648 1820 77654
rect 1768 77590 1820 77596
rect 1676 77376 1728 77382
rect 1676 77318 1728 77324
rect 1492 77036 1544 77042
rect 1492 76978 1544 76984
rect 1398 76936 1454 76945
rect 1398 76871 1454 76880
rect 1584 76832 1636 76838
rect 1584 76774 1636 76780
rect 1400 76424 1452 76430
rect 1306 76392 1362 76401
rect 1400 76366 1452 76372
rect 1306 76327 1362 76336
rect 1308 75948 1360 75954
rect 1308 75890 1360 75896
rect 1320 74769 1348 75890
rect 1412 75857 1440 76366
rect 1492 76288 1544 76294
rect 1492 76230 1544 76236
rect 1398 75848 1454 75857
rect 1398 75783 1454 75792
rect 1400 75336 1452 75342
rect 1400 75278 1452 75284
rect 1306 74760 1362 74769
rect 1124 74724 1176 74730
rect 1306 74695 1362 74704
rect 1124 74666 1176 74672
rect 480 73568 532 73574
rect 480 73510 532 73516
rect 204 52964 256 52970
rect 204 52906 256 52912
rect 112 46504 164 46510
rect 112 46446 164 46452
rect 20 45008 72 45014
rect 20 44950 72 44956
rect 32 36582 60 44950
rect 20 36576 72 36582
rect 20 36518 72 36524
rect 124 27470 152 46446
rect 216 35222 244 52906
rect 296 39364 348 39370
rect 296 39306 348 39312
rect 204 35216 256 35222
rect 204 35158 256 35164
rect 204 31748 256 31754
rect 204 31690 256 31696
rect 112 27464 164 27470
rect 112 27406 164 27412
rect 216 12442 244 31690
rect 308 19446 336 39306
rect 388 37392 440 37398
rect 388 37334 440 37340
rect 296 19440 348 19446
rect 296 19382 348 19388
rect 400 18154 428 37334
rect 492 36378 520 73510
rect 848 73024 900 73030
rect 848 72966 900 72972
rect 756 66088 808 66094
rect 756 66030 808 66036
rect 768 60734 796 66030
rect 860 65210 888 72966
rect 1136 65736 1164 74666
rect 1412 73681 1440 75278
rect 1504 73846 1532 76230
rect 1596 74322 1624 76774
rect 1688 74934 1716 77318
rect 1676 74928 1728 74934
rect 1676 74870 1728 74876
rect 1676 74792 1728 74798
rect 1676 74734 1728 74740
rect 1584 74316 1636 74322
rect 1584 74258 1636 74264
rect 1584 74180 1636 74186
rect 1584 74122 1636 74128
rect 1492 73840 1544 73846
rect 1492 73782 1544 73788
rect 1398 73672 1454 73681
rect 1398 73607 1454 73616
rect 1492 73636 1544 73642
rect 1492 73578 1544 73584
rect 1504 73166 1532 73578
rect 1596 73370 1624 74122
rect 1688 74118 1716 74734
rect 1676 74112 1728 74118
rect 1676 74054 1728 74060
rect 1688 73642 1716 74054
rect 1676 73636 1728 73642
rect 1676 73578 1728 73584
rect 1584 73364 1636 73370
rect 1584 73306 1636 73312
rect 1492 73160 1544 73166
rect 1492 73102 1544 73108
rect 1676 73160 1728 73166
rect 1780 73148 1808 77590
rect 2976 77518 3004 77959
rect 2044 77512 2096 77518
rect 2042 77480 2044 77489
rect 2964 77512 3016 77518
rect 2096 77480 2098 77489
rect 2964 77454 3016 77460
rect 2042 77415 2098 77424
rect 2504 77376 2556 77382
rect 2504 77318 2556 77324
rect 2228 76832 2280 76838
rect 2228 76774 2280 76780
rect 2044 75336 2096 75342
rect 2042 75304 2044 75313
rect 2096 75304 2098 75313
rect 2042 75239 2098 75248
rect 2240 74934 2268 76774
rect 2228 74928 2280 74934
rect 2228 74870 2280 74876
rect 2136 74860 2188 74866
rect 2136 74802 2188 74808
rect 2148 74254 2176 74802
rect 2516 74338 2544 77318
rect 3068 77042 3096 79047
rect 3804 77518 3832 79591
rect 9586 79520 9642 79529
rect 9586 79455 9642 79464
rect 9494 78024 9550 78033
rect 9494 77959 9550 77968
rect 5845 77820 6153 77840
rect 5845 77818 5851 77820
rect 5907 77818 5931 77820
rect 5987 77818 6011 77820
rect 6067 77818 6091 77820
rect 6147 77818 6153 77820
rect 5907 77766 5909 77818
rect 6089 77766 6091 77818
rect 5845 77764 5851 77766
rect 5907 77764 5931 77766
rect 5987 77764 6011 77766
rect 6067 77764 6091 77766
rect 6147 77764 6153 77766
rect 5845 77744 6153 77764
rect 9109 77820 9417 77840
rect 9109 77818 9115 77820
rect 9171 77818 9195 77820
rect 9251 77818 9275 77820
rect 9331 77818 9355 77820
rect 9411 77818 9417 77820
rect 9171 77766 9173 77818
rect 9353 77766 9355 77818
rect 9109 77764 9115 77766
rect 9171 77764 9195 77766
rect 9251 77764 9275 77766
rect 9331 77764 9355 77766
rect 9411 77764 9417 77766
rect 9109 77744 9417 77764
rect 9508 77722 9536 77959
rect 9496 77716 9548 77722
rect 9496 77658 9548 77664
rect 3792 77512 3844 77518
rect 3792 77454 3844 77460
rect 5540 77512 5592 77518
rect 5540 77454 5592 77460
rect 3976 77376 4028 77382
rect 3976 77318 4028 77324
rect 3056 77036 3108 77042
rect 3056 76978 3108 76984
rect 3608 76832 3660 76838
rect 3608 76774 3660 76780
rect 2582 76732 2890 76752
rect 2582 76730 2588 76732
rect 2644 76730 2668 76732
rect 2724 76730 2748 76732
rect 2804 76730 2828 76732
rect 2884 76730 2890 76732
rect 2644 76678 2646 76730
rect 2826 76678 2828 76730
rect 2582 76676 2588 76678
rect 2644 76676 2668 76678
rect 2724 76676 2748 76678
rect 2804 76676 2828 76678
rect 2884 76676 2890 76678
rect 2582 76656 2890 76676
rect 3056 76084 3108 76090
rect 3056 76026 3108 76032
rect 2582 75644 2890 75664
rect 2582 75642 2588 75644
rect 2644 75642 2668 75644
rect 2724 75642 2748 75644
rect 2804 75642 2828 75644
rect 2884 75642 2890 75644
rect 2644 75590 2646 75642
rect 2826 75590 2828 75642
rect 2582 75588 2588 75590
rect 2644 75588 2668 75590
rect 2724 75588 2748 75590
rect 2804 75588 2828 75590
rect 2884 75588 2890 75590
rect 2582 75568 2890 75588
rect 2964 75200 3016 75206
rect 2964 75142 3016 75148
rect 2596 74860 2648 74866
rect 2596 74802 2648 74808
rect 2608 74730 2636 74802
rect 2596 74724 2648 74730
rect 2596 74666 2648 74672
rect 2582 74556 2890 74576
rect 2582 74554 2588 74556
rect 2644 74554 2668 74556
rect 2724 74554 2748 74556
rect 2804 74554 2828 74556
rect 2884 74554 2890 74556
rect 2644 74502 2646 74554
rect 2826 74502 2828 74554
rect 2582 74500 2588 74502
rect 2644 74500 2668 74502
rect 2724 74500 2748 74502
rect 2804 74500 2828 74502
rect 2884 74500 2890 74502
rect 2582 74480 2890 74500
rect 2516 74310 2728 74338
rect 2700 74254 2728 74310
rect 2136 74248 2188 74254
rect 2136 74190 2188 74196
rect 2688 74248 2740 74254
rect 2688 74190 2740 74196
rect 2780 74248 2832 74254
rect 2780 74190 2832 74196
rect 2148 73778 2176 74190
rect 2504 74112 2556 74118
rect 2504 74054 2556 74060
rect 2516 73914 2544 74054
rect 2504 73908 2556 73914
rect 2504 73850 2556 73856
rect 2136 73772 2188 73778
rect 2136 73714 2188 73720
rect 2412 73772 2464 73778
rect 2412 73714 2464 73720
rect 2148 73166 2176 73714
rect 2424 73166 2452 73714
rect 2792 73710 2820 74190
rect 2976 73846 3004 75142
rect 2964 73840 3016 73846
rect 2964 73782 3016 73788
rect 2780 73704 2832 73710
rect 2780 73646 2832 73652
rect 2964 73704 3016 73710
rect 2964 73646 3016 73652
rect 2582 73468 2890 73488
rect 2582 73466 2588 73468
rect 2644 73466 2668 73468
rect 2724 73466 2748 73468
rect 2804 73466 2828 73468
rect 2884 73466 2890 73468
rect 2644 73414 2646 73466
rect 2826 73414 2828 73466
rect 2582 73412 2588 73414
rect 2644 73412 2668 73414
rect 2724 73412 2748 73414
rect 2804 73412 2828 73414
rect 2884 73412 2890 73414
rect 2582 73392 2890 73412
rect 2976 73250 3004 73646
rect 2884 73222 3004 73250
rect 2884 73166 2912 73222
rect 1728 73120 1808 73148
rect 2136 73160 2188 73166
rect 1676 73102 1728 73108
rect 2136 73102 2188 73108
rect 2412 73160 2464 73166
rect 2412 73102 2464 73108
rect 2872 73160 2924 73166
rect 2872 73102 2924 73108
rect 2964 73160 3016 73166
rect 3068 73148 3096 76026
rect 3148 75472 3200 75478
rect 3148 75414 3200 75420
rect 3016 73120 3096 73148
rect 2964 73102 3016 73108
rect 1504 72758 1532 73102
rect 1584 73092 1636 73098
rect 1584 73034 1636 73040
rect 1492 72752 1544 72758
rect 1492 72694 1544 72700
rect 1400 72684 1452 72690
rect 1400 72626 1452 72632
rect 1412 72457 1440 72626
rect 1596 72622 1624 73034
rect 2042 72992 2098 73001
rect 2042 72927 2098 72936
rect 2056 72690 2084 72927
rect 2148 72690 2176 73102
rect 2044 72684 2096 72690
rect 2044 72626 2096 72632
rect 2136 72684 2188 72690
rect 2136 72626 2188 72632
rect 1584 72616 1636 72622
rect 1584 72558 1636 72564
rect 1676 72480 1728 72486
rect 1398 72448 1454 72457
rect 1676 72422 1728 72428
rect 2320 72480 2372 72486
rect 2320 72422 2372 72428
rect 1398 72383 1454 72392
rect 1400 72072 1452 72078
rect 1400 72014 1452 72020
rect 1412 71913 1440 72014
rect 1398 71904 1454 71913
rect 1398 71839 1454 71848
rect 1400 71596 1452 71602
rect 1400 71538 1452 71544
rect 1412 71369 1440 71538
rect 1398 71360 1454 71369
rect 1398 71295 1454 71304
rect 1400 70984 1452 70990
rect 1400 70926 1452 70932
rect 1412 70825 1440 70926
rect 1398 70816 1454 70825
rect 1398 70751 1454 70760
rect 1400 70508 1452 70514
rect 1400 70450 1452 70456
rect 1412 70281 1440 70450
rect 1398 70272 1454 70281
rect 1398 70207 1454 70216
rect 1400 69896 1452 69902
rect 1400 69838 1452 69844
rect 1412 69737 1440 69838
rect 1398 69728 1454 69737
rect 1398 69663 1454 69672
rect 1400 69420 1452 69426
rect 1400 69362 1452 69368
rect 1412 69193 1440 69362
rect 1398 69184 1454 69193
rect 1398 69119 1454 69128
rect 1400 68808 1452 68814
rect 1400 68750 1452 68756
rect 1412 68649 1440 68750
rect 1492 68672 1544 68678
rect 1398 68640 1454 68649
rect 1492 68614 1544 68620
rect 1398 68575 1454 68584
rect 1400 68332 1452 68338
rect 1400 68274 1452 68280
rect 1412 68105 1440 68274
rect 1398 68096 1454 68105
rect 1398 68031 1454 68040
rect 1400 67720 1452 67726
rect 1400 67662 1452 67668
rect 1216 67244 1268 67250
rect 1216 67186 1268 67192
rect 1228 65793 1256 67186
rect 1308 66632 1360 66638
rect 1308 66574 1360 66580
rect 1044 65708 1164 65736
rect 1214 65784 1270 65793
rect 1214 65719 1270 65728
rect 1044 65498 1072 65708
rect 1044 65470 1164 65498
rect 1032 65408 1084 65414
rect 1032 65350 1084 65356
rect 848 65204 900 65210
rect 848 65146 900 65152
rect 768 60706 980 60734
rect 848 53168 900 53174
rect 848 53110 900 53116
rect 756 52624 808 52630
rect 756 52566 808 52572
rect 664 49292 716 49298
rect 664 49234 716 49240
rect 572 48680 624 48686
rect 572 48622 624 48628
rect 480 36372 532 36378
rect 480 36314 532 36320
rect 480 35624 532 35630
rect 480 35566 532 35572
rect 388 18148 440 18154
rect 388 18090 440 18096
rect 492 13802 520 35566
rect 584 21690 612 48622
rect 676 27538 704 49234
rect 768 47666 796 52566
rect 756 47660 808 47666
rect 756 47602 808 47608
rect 860 47546 888 53110
rect 768 47518 888 47546
rect 768 38214 796 47518
rect 848 47456 900 47462
rect 848 47398 900 47404
rect 756 38208 808 38214
rect 756 38150 808 38156
rect 756 36576 808 36582
rect 756 36518 808 36524
rect 664 27532 716 27538
rect 664 27474 716 27480
rect 572 21684 624 21690
rect 572 21626 624 21632
rect 768 20874 796 36518
rect 860 28966 888 47398
rect 952 33114 980 60706
rect 940 33108 992 33114
rect 940 33050 992 33056
rect 1044 32570 1072 65350
rect 1136 39098 1164 65470
rect 1320 65249 1348 66574
rect 1412 66337 1440 67662
rect 1398 66328 1454 66337
rect 1398 66263 1454 66272
rect 1400 65544 1452 65550
rect 1400 65486 1452 65492
rect 1306 65240 1362 65249
rect 1216 65204 1268 65210
rect 1306 65175 1362 65184
rect 1216 65146 1268 65152
rect 1124 39092 1176 39098
rect 1124 39034 1176 39040
rect 1124 36712 1176 36718
rect 1124 36654 1176 36660
rect 1032 32564 1084 32570
rect 1032 32506 1084 32512
rect 940 30864 992 30870
rect 940 30806 992 30812
rect 848 28960 900 28966
rect 848 28902 900 28908
rect 952 28778 980 30806
rect 860 28750 980 28778
rect 860 26234 888 28750
rect 1032 28416 1084 28422
rect 1032 28358 1084 28364
rect 940 28144 992 28150
rect 940 28086 992 28092
rect 952 27062 980 28086
rect 940 27056 992 27062
rect 940 26998 992 27004
rect 860 26206 980 26234
rect 756 20868 808 20874
rect 756 20810 808 20816
rect 480 13796 532 13802
rect 480 13738 532 13744
rect 204 12436 256 12442
rect 204 12378 256 12384
rect 952 9110 980 26206
rect 940 9104 992 9110
rect 940 9046 992 9052
rect 1044 5778 1072 28358
rect 1136 12782 1164 36654
rect 1228 35290 1256 65146
rect 1308 65068 1360 65074
rect 1308 65010 1360 65016
rect 1320 63617 1348 65010
rect 1412 64705 1440 65486
rect 1398 64696 1454 64705
rect 1398 64631 1454 64640
rect 1400 64456 1452 64462
rect 1400 64398 1452 64404
rect 1412 64002 1440 64398
rect 1504 64122 1532 68614
rect 1584 67040 1636 67046
rect 1584 66982 1636 66988
rect 1492 64116 1544 64122
rect 1492 64058 1544 64064
rect 1490 64016 1546 64025
rect 1412 63974 1490 64002
rect 1490 63951 1492 63960
rect 1544 63951 1546 63960
rect 1492 63922 1544 63928
rect 1306 63608 1362 63617
rect 1306 63543 1362 63552
rect 1504 63374 1532 63922
rect 1492 63368 1544 63374
rect 1492 63310 1544 63316
rect 1504 62898 1532 63310
rect 1492 62892 1544 62898
rect 1492 62834 1544 62840
rect 1492 62144 1544 62150
rect 1492 62086 1544 62092
rect 1400 61600 1452 61606
rect 1400 61542 1452 61548
rect 1412 60897 1440 61542
rect 1504 61441 1532 62086
rect 1490 61432 1546 61441
rect 1490 61367 1546 61376
rect 1492 61056 1544 61062
rect 1492 60998 1544 61004
rect 1398 60888 1454 60897
rect 1398 60823 1454 60832
rect 1400 60512 1452 60518
rect 1400 60454 1452 60460
rect 1412 59673 1440 60454
rect 1504 60353 1532 60998
rect 1490 60344 1546 60353
rect 1490 60279 1546 60288
rect 1492 59968 1544 59974
rect 1492 59910 1544 59916
rect 1398 59664 1454 59673
rect 1398 59599 1454 59608
rect 1400 59424 1452 59430
rect 1400 59366 1452 59372
rect 1412 58585 1440 59366
rect 1504 59129 1532 59910
rect 1490 59120 1546 59129
rect 1490 59055 1546 59064
rect 1492 58880 1544 58886
rect 1492 58822 1544 58828
rect 1398 58576 1454 58585
rect 1398 58511 1454 58520
rect 1400 58336 1452 58342
rect 1400 58278 1452 58284
rect 1308 58064 1360 58070
rect 1308 58006 1360 58012
rect 1320 52698 1348 58006
rect 1412 56953 1440 58278
rect 1504 58041 1532 58822
rect 1490 58032 1546 58041
rect 1490 57967 1546 57976
rect 1492 57928 1544 57934
rect 1596 57882 1624 66982
rect 1688 66230 1716 72422
rect 2332 71670 2360 72422
rect 2424 72078 2452 73102
rect 2504 72480 2556 72486
rect 2884 72468 2912 73102
rect 2884 72440 3004 72468
rect 2504 72422 2556 72428
rect 2516 72214 2544 72422
rect 2582 72380 2890 72400
rect 2582 72378 2588 72380
rect 2644 72378 2668 72380
rect 2724 72378 2748 72380
rect 2804 72378 2828 72380
rect 2884 72378 2890 72380
rect 2644 72326 2646 72378
rect 2826 72326 2828 72378
rect 2582 72324 2588 72326
rect 2644 72324 2668 72326
rect 2724 72324 2748 72326
rect 2804 72324 2828 72326
rect 2884 72324 2890 72326
rect 2582 72304 2890 72324
rect 2504 72208 2556 72214
rect 2504 72150 2556 72156
rect 2976 72078 3004 72440
rect 3160 72146 3188 75414
rect 3516 74792 3568 74798
rect 3516 74734 3568 74740
rect 3332 74180 3384 74186
rect 3332 74122 3384 74128
rect 3148 72140 3200 72146
rect 3148 72082 3200 72088
rect 2412 72072 2464 72078
rect 2412 72014 2464 72020
rect 2964 72072 3016 72078
rect 2964 72014 3016 72020
rect 2872 71936 2924 71942
rect 2872 71878 2924 71884
rect 2320 71664 2372 71670
rect 2320 71606 2372 71612
rect 2884 71534 2912 71878
rect 2976 71602 3004 72014
rect 2964 71596 3016 71602
rect 2964 71538 3016 71544
rect 2872 71528 2924 71534
rect 2872 71470 2924 71476
rect 2504 71392 2556 71398
rect 2504 71334 2556 71340
rect 2412 70848 2464 70854
rect 2412 70790 2464 70796
rect 2044 70644 2096 70650
rect 2044 70586 2096 70592
rect 1768 69216 1820 69222
rect 1768 69158 1820 69164
rect 1676 66224 1728 66230
rect 1676 66166 1728 66172
rect 1676 65408 1728 65414
rect 1676 65350 1728 65356
rect 1544 57876 1624 57882
rect 1492 57870 1624 57876
rect 1504 57854 1624 57870
rect 1492 57792 1544 57798
rect 1492 57734 1544 57740
rect 1582 57760 1638 57769
rect 1504 57458 1532 57734
rect 1582 57695 1638 57704
rect 1492 57452 1544 57458
rect 1492 57394 1544 57400
rect 1398 56944 1454 56953
rect 1398 56879 1454 56888
rect 1400 56840 1452 56846
rect 1504 56828 1532 57394
rect 1452 56800 1532 56828
rect 1400 56782 1452 56788
rect 1412 56370 1440 56782
rect 1400 56364 1452 56370
rect 1452 56324 1532 56352
rect 1400 56306 1452 56312
rect 1400 55820 1452 55826
rect 1504 55808 1532 56324
rect 1452 55780 1532 55808
rect 1400 55762 1452 55768
rect 1412 55282 1440 55762
rect 1400 55276 1452 55282
rect 1400 55218 1452 55224
rect 1596 55214 1624 57695
rect 1688 57526 1716 65350
rect 1780 64462 1808 69158
rect 1860 68128 1912 68134
rect 1860 68070 1912 68076
rect 1768 64456 1820 64462
rect 1768 64398 1820 64404
rect 1768 63572 1820 63578
rect 1768 63514 1820 63520
rect 1780 63186 1808 63514
rect 1872 63374 1900 68070
rect 1952 67856 2004 67862
rect 1952 67798 2004 67804
rect 1860 63368 1912 63374
rect 1860 63310 1912 63316
rect 1780 63158 1900 63186
rect 1768 62892 1820 62898
rect 1768 62834 1820 62840
rect 1780 62354 1808 62834
rect 1768 62348 1820 62354
rect 1768 62290 1820 62296
rect 1768 61600 1820 61606
rect 1768 61542 1820 61548
rect 1780 59158 1808 61542
rect 1768 59152 1820 59158
rect 1768 59094 1820 59100
rect 1768 59016 1820 59022
rect 1768 58958 1820 58964
rect 1676 57520 1728 57526
rect 1676 57462 1728 57468
rect 1676 56500 1728 56506
rect 1676 56442 1728 56448
rect 1688 55282 1716 56442
rect 1676 55276 1728 55282
rect 1676 55218 1728 55224
rect 1584 55208 1636 55214
rect 1584 55150 1636 55156
rect 1400 55140 1452 55146
rect 1400 55082 1452 55088
rect 1412 54754 1440 55082
rect 1412 54726 1624 54754
rect 1400 54664 1452 54670
rect 1400 54606 1452 54612
rect 1308 52692 1360 52698
rect 1308 52634 1360 52640
rect 1412 51074 1440 54606
rect 1492 54528 1544 54534
rect 1492 54470 1544 54476
rect 1504 54233 1532 54470
rect 1490 54224 1546 54233
rect 1490 54159 1546 54168
rect 1492 53984 1544 53990
rect 1492 53926 1544 53932
rect 1504 53689 1532 53926
rect 1490 53680 1546 53689
rect 1490 53615 1546 53624
rect 1492 53236 1544 53242
rect 1492 53178 1544 53184
rect 1504 53009 1532 53178
rect 1490 53000 1546 53009
rect 1490 52935 1546 52944
rect 1492 52896 1544 52902
rect 1492 52838 1544 52844
rect 1504 52465 1532 52838
rect 1490 52456 1546 52465
rect 1490 52391 1546 52400
rect 1492 52352 1544 52358
rect 1492 52294 1544 52300
rect 1504 51377 1532 52294
rect 1490 51368 1546 51377
rect 1490 51303 1546 51312
rect 1596 51270 1624 54726
rect 1676 52692 1728 52698
rect 1676 52634 1728 52640
rect 1688 51406 1716 52634
rect 1676 51400 1728 51406
rect 1676 51342 1728 51348
rect 1492 51264 1544 51270
rect 1492 51206 1544 51212
rect 1584 51264 1636 51270
rect 1584 51206 1636 51212
rect 1320 51046 1440 51074
rect 1320 50130 1348 51046
rect 1400 50924 1452 50930
rect 1400 50866 1452 50872
rect 1412 50318 1440 50866
rect 1504 50318 1532 51206
rect 1676 50992 1728 50998
rect 1674 50960 1676 50969
rect 1728 50960 1730 50969
rect 1674 50895 1730 50904
rect 1400 50312 1452 50318
rect 1400 50254 1452 50260
rect 1492 50312 1544 50318
rect 1492 50254 1544 50260
rect 1320 50102 1440 50130
rect 1412 45554 1440 50102
rect 1780 49978 1808 58958
rect 1872 56710 1900 63158
rect 1964 62898 1992 67798
rect 2056 65142 2084 70586
rect 2320 69760 2372 69766
rect 2320 69702 2372 69708
rect 2136 67924 2188 67930
rect 2136 67866 2188 67872
rect 2044 65136 2096 65142
rect 2044 65078 2096 65084
rect 2148 63594 2176 67866
rect 2228 67720 2280 67726
rect 2228 67662 2280 67668
rect 2240 67561 2268 67662
rect 2226 67552 2282 67561
rect 2226 67487 2282 67496
rect 2228 67244 2280 67250
rect 2228 67186 2280 67192
rect 2240 67017 2268 67186
rect 2332 67182 2360 69702
rect 2320 67176 2372 67182
rect 2320 67118 2372 67124
rect 2320 67040 2372 67046
rect 2226 67008 2282 67017
rect 2320 66982 2372 66988
rect 2226 66943 2282 66952
rect 2228 66632 2280 66638
rect 2228 66574 2280 66580
rect 2240 66298 2268 66574
rect 2228 66292 2280 66298
rect 2228 66234 2280 66240
rect 2240 65618 2268 66234
rect 2228 65612 2280 65618
rect 2228 65554 2280 65560
rect 2240 65074 2268 65554
rect 2228 65068 2280 65074
rect 2228 65010 2280 65016
rect 2228 64932 2280 64938
rect 2228 64874 2280 64880
rect 2056 63578 2176 63594
rect 2044 63572 2176 63578
rect 2096 63566 2176 63572
rect 2044 63514 2096 63520
rect 2044 63368 2096 63374
rect 2044 63310 2096 63316
rect 2056 62898 2084 63310
rect 1952 62892 2004 62898
rect 1952 62834 2004 62840
rect 2044 62892 2096 62898
rect 2044 62834 2096 62840
rect 2240 62778 2268 64874
rect 2332 63578 2360 66982
rect 2424 66774 2452 70790
rect 2412 66768 2464 66774
rect 2412 66710 2464 66716
rect 2516 66638 2544 71334
rect 2582 71292 2890 71312
rect 2582 71290 2588 71292
rect 2644 71290 2668 71292
rect 2724 71290 2748 71292
rect 2804 71290 2828 71292
rect 2884 71290 2890 71292
rect 2644 71238 2646 71290
rect 2826 71238 2828 71290
rect 2582 71236 2588 71238
rect 2644 71236 2668 71238
rect 2724 71236 2748 71238
rect 2804 71236 2828 71238
rect 2884 71236 2890 71238
rect 2582 71216 2890 71236
rect 2582 70204 2890 70224
rect 2582 70202 2588 70204
rect 2644 70202 2668 70204
rect 2724 70202 2748 70204
rect 2804 70202 2828 70204
rect 2884 70202 2890 70204
rect 2644 70150 2646 70202
rect 2826 70150 2828 70202
rect 2582 70148 2588 70150
rect 2644 70148 2668 70150
rect 2724 70148 2748 70150
rect 2804 70148 2828 70150
rect 2884 70148 2890 70150
rect 2582 70128 2890 70148
rect 2582 69116 2890 69136
rect 2582 69114 2588 69116
rect 2644 69114 2668 69116
rect 2724 69114 2748 69116
rect 2804 69114 2828 69116
rect 2884 69114 2890 69116
rect 2644 69062 2646 69114
rect 2826 69062 2828 69114
rect 2582 69060 2588 69062
rect 2644 69060 2668 69062
rect 2724 69060 2748 69062
rect 2804 69060 2828 69062
rect 2884 69060 2890 69062
rect 2582 69040 2890 69060
rect 3344 69018 3372 74122
rect 3528 73778 3556 74734
rect 3620 73846 3648 76774
rect 3700 74860 3752 74866
rect 3700 74802 3752 74808
rect 3712 74186 3740 74802
rect 3988 74254 4016 77318
rect 4213 77276 4521 77296
rect 4213 77274 4219 77276
rect 4275 77274 4299 77276
rect 4355 77274 4379 77276
rect 4435 77274 4459 77276
rect 4515 77274 4521 77276
rect 4275 77222 4277 77274
rect 4457 77222 4459 77274
rect 4213 77220 4219 77222
rect 4275 77220 4299 77222
rect 4355 77220 4379 77222
rect 4435 77220 4459 77222
rect 4515 77220 4521 77222
rect 4213 77200 4521 77220
rect 4213 76188 4521 76208
rect 4213 76186 4219 76188
rect 4275 76186 4299 76188
rect 4355 76186 4379 76188
rect 4435 76186 4459 76188
rect 4515 76186 4521 76188
rect 4275 76134 4277 76186
rect 4457 76134 4459 76186
rect 4213 76132 4219 76134
rect 4275 76132 4299 76134
rect 4355 76132 4379 76134
rect 4435 76132 4459 76134
rect 4515 76132 4521 76134
rect 4213 76112 4521 76132
rect 4213 75100 4521 75120
rect 4213 75098 4219 75100
rect 4275 75098 4299 75100
rect 4355 75098 4379 75100
rect 4435 75098 4459 75100
rect 4515 75098 4521 75100
rect 4275 75046 4277 75098
rect 4457 75046 4459 75098
rect 4213 75044 4219 75046
rect 4275 75044 4299 75046
rect 4355 75044 4379 75046
rect 4435 75044 4459 75046
rect 4515 75044 4521 75046
rect 4213 75024 4521 75044
rect 5552 75002 5580 77454
rect 7477 77276 7785 77296
rect 7477 77274 7483 77276
rect 7539 77274 7563 77276
rect 7619 77274 7643 77276
rect 7699 77274 7723 77276
rect 7779 77274 7785 77276
rect 7539 77222 7541 77274
rect 7721 77222 7723 77274
rect 7477 77220 7483 77222
rect 7539 77220 7563 77222
rect 7619 77220 7643 77222
rect 7699 77220 7723 77222
rect 7779 77220 7785 77222
rect 7477 77200 7785 77220
rect 9600 77178 9628 79455
rect 10966 78704 11022 78713
rect 10966 78639 10968 78648
rect 11020 78639 11022 78648
rect 10968 78610 11020 78616
rect 10048 77376 10100 77382
rect 10048 77318 10100 77324
rect 10060 77217 10088 77318
rect 10046 77208 10102 77217
rect 9588 77172 9640 77178
rect 10046 77143 10102 77152
rect 9588 77114 9640 77120
rect 8300 77036 8352 77042
rect 8300 76978 8352 76984
rect 9680 77036 9732 77042
rect 9680 76978 9732 76984
rect 5845 76732 6153 76752
rect 5845 76730 5851 76732
rect 5907 76730 5931 76732
rect 5987 76730 6011 76732
rect 6067 76730 6091 76732
rect 6147 76730 6153 76732
rect 5907 76678 5909 76730
rect 6089 76678 6091 76730
rect 5845 76676 5851 76678
rect 5907 76676 5931 76678
rect 5987 76676 6011 76678
rect 6067 76676 6091 76678
rect 6147 76676 6153 76678
rect 5845 76656 6153 76676
rect 7477 76188 7785 76208
rect 7477 76186 7483 76188
rect 7539 76186 7563 76188
rect 7619 76186 7643 76188
rect 7699 76186 7723 76188
rect 7779 76186 7785 76188
rect 7539 76134 7541 76186
rect 7721 76134 7723 76186
rect 7477 76132 7483 76134
rect 7539 76132 7563 76134
rect 7619 76132 7643 76134
rect 7699 76132 7723 76134
rect 7779 76132 7785 76134
rect 7477 76112 7785 76132
rect 6276 75880 6328 75886
rect 6276 75822 6328 75828
rect 5845 75644 6153 75664
rect 5845 75642 5851 75644
rect 5907 75642 5931 75644
rect 5987 75642 6011 75644
rect 6067 75642 6091 75644
rect 6147 75642 6153 75644
rect 5907 75590 5909 75642
rect 6089 75590 6091 75642
rect 5845 75588 5851 75590
rect 5907 75588 5931 75590
rect 5987 75588 6011 75590
rect 6067 75588 6091 75590
rect 6147 75588 6153 75590
rect 5845 75568 6153 75588
rect 5540 74996 5592 75002
rect 5540 74938 5592 74944
rect 6288 74662 6316 75822
rect 7477 75100 7785 75120
rect 7477 75098 7483 75100
rect 7539 75098 7563 75100
rect 7619 75098 7643 75100
rect 7699 75098 7723 75100
rect 7779 75098 7785 75100
rect 7539 75046 7541 75098
rect 7721 75046 7723 75098
rect 7477 75044 7483 75046
rect 7539 75044 7563 75046
rect 7619 75044 7643 75046
rect 7699 75044 7723 75046
rect 7779 75044 7785 75046
rect 7477 75024 7785 75044
rect 6552 74928 6604 74934
rect 6552 74870 6604 74876
rect 6276 74656 6328 74662
rect 6276 74598 6328 74604
rect 5845 74556 6153 74576
rect 5845 74554 5851 74556
rect 5907 74554 5931 74556
rect 5987 74554 6011 74556
rect 6067 74554 6091 74556
rect 6147 74554 6153 74556
rect 5907 74502 5909 74554
rect 6089 74502 6091 74554
rect 5845 74500 5851 74502
rect 5907 74500 5931 74502
rect 5987 74500 6011 74502
rect 6067 74500 6091 74502
rect 6147 74500 6153 74502
rect 5845 74480 6153 74500
rect 5632 74316 5684 74322
rect 5632 74258 5684 74264
rect 3792 74248 3844 74254
rect 3790 74216 3792 74225
rect 3976 74248 4028 74254
rect 3844 74216 3846 74225
rect 3700 74180 3752 74186
rect 3976 74190 4028 74196
rect 4804 74248 4856 74254
rect 4804 74190 4856 74196
rect 3790 74151 3846 74160
rect 3700 74122 3752 74128
rect 3608 73840 3660 73846
rect 3608 73782 3660 73788
rect 3516 73772 3568 73778
rect 3516 73714 3568 73720
rect 3528 73234 3556 73714
rect 3712 73658 3740 74122
rect 4068 74112 4120 74118
rect 4068 74054 4120 74060
rect 3792 73704 3844 73710
rect 3712 73652 3792 73658
rect 3712 73646 3844 73652
rect 3712 73630 3832 73646
rect 3516 73228 3568 73234
rect 3516 73170 3568 73176
rect 3332 69012 3384 69018
rect 3332 68954 3384 68960
rect 2582 68028 2890 68048
rect 2582 68026 2588 68028
rect 2644 68026 2668 68028
rect 2724 68026 2748 68028
rect 2804 68026 2828 68028
rect 2884 68026 2890 68028
rect 2644 67974 2646 68026
rect 2826 67974 2828 68026
rect 2582 67972 2588 67974
rect 2644 67972 2668 67974
rect 2724 67972 2748 67974
rect 2804 67972 2828 67974
rect 2884 67972 2890 67974
rect 2582 67952 2890 67972
rect 3056 67176 3108 67182
rect 3056 67118 3108 67124
rect 2582 66940 2890 66960
rect 2582 66938 2588 66940
rect 2644 66938 2668 66940
rect 2724 66938 2748 66940
rect 2804 66938 2828 66940
rect 2884 66938 2890 66940
rect 2644 66886 2646 66938
rect 2826 66886 2828 66938
rect 2582 66884 2588 66886
rect 2644 66884 2668 66886
rect 2724 66884 2748 66886
rect 2804 66884 2828 66886
rect 2884 66884 2890 66886
rect 2582 66864 2890 66884
rect 2688 66768 2740 66774
rect 2688 66710 2740 66716
rect 2504 66632 2556 66638
rect 2504 66574 2556 66580
rect 2412 66496 2464 66502
rect 2412 66438 2464 66444
rect 2320 63572 2372 63578
rect 2320 63514 2372 63520
rect 1952 62756 2004 62762
rect 1952 62698 2004 62704
rect 2044 62756 2096 62762
rect 2240 62750 2360 62778
rect 2044 62698 2096 62704
rect 1964 62150 1992 62698
rect 2056 62642 2084 62698
rect 2056 62614 2268 62642
rect 2044 62484 2096 62490
rect 2044 62426 2096 62432
rect 1952 62144 2004 62150
rect 1952 62086 2004 62092
rect 1952 58540 2004 58546
rect 1952 58482 2004 58488
rect 1964 57905 1992 58482
rect 1950 57896 2006 57905
rect 1950 57831 2006 57840
rect 1952 57792 2004 57798
rect 1952 57734 2004 57740
rect 1964 57594 1992 57734
rect 1952 57588 2004 57594
rect 1952 57530 2004 57536
rect 1952 57452 2004 57458
rect 1952 57394 2004 57400
rect 1964 56846 1992 57394
rect 1952 56840 2004 56846
rect 1952 56782 2004 56788
rect 2056 56778 2084 62426
rect 2136 62144 2188 62150
rect 2136 62086 2188 62092
rect 2148 59242 2176 62086
rect 2240 59401 2268 62614
rect 2332 62370 2360 62750
rect 2424 62490 2452 66438
rect 2700 66162 2728 66710
rect 2872 66632 2924 66638
rect 2872 66574 2924 66580
rect 2884 66298 2912 66574
rect 2872 66292 2924 66298
rect 2872 66234 2924 66240
rect 2884 66162 2912 66234
rect 2504 66156 2556 66162
rect 2504 66098 2556 66104
rect 2688 66156 2740 66162
rect 2688 66098 2740 66104
rect 2872 66156 2924 66162
rect 2924 66116 3004 66144
rect 2872 66098 2924 66104
rect 2516 65006 2544 66098
rect 2582 65852 2890 65872
rect 2582 65850 2588 65852
rect 2644 65850 2668 65852
rect 2724 65850 2748 65852
rect 2804 65850 2828 65852
rect 2884 65850 2890 65852
rect 2644 65798 2646 65850
rect 2826 65798 2828 65850
rect 2582 65796 2588 65798
rect 2644 65796 2668 65798
rect 2724 65796 2748 65798
rect 2804 65796 2828 65798
rect 2884 65796 2890 65798
rect 2582 65776 2890 65796
rect 2976 65074 3004 66116
rect 2964 65068 3016 65074
rect 2964 65010 3016 65016
rect 2504 65000 2556 65006
rect 2504 64942 2556 64948
rect 2582 64764 2890 64784
rect 2582 64762 2588 64764
rect 2644 64762 2668 64764
rect 2724 64762 2748 64764
rect 2804 64762 2828 64764
rect 2884 64762 2890 64764
rect 2644 64710 2646 64762
rect 2826 64710 2828 64762
rect 2582 64708 2588 64710
rect 2644 64708 2668 64710
rect 2724 64708 2748 64710
rect 2804 64708 2828 64710
rect 2884 64708 2890 64710
rect 2582 64688 2890 64708
rect 2964 64524 3016 64530
rect 2964 64466 3016 64472
rect 2780 64456 2832 64462
rect 2780 64398 2832 64404
rect 2872 64456 2924 64462
rect 2872 64398 2924 64404
rect 2792 64161 2820 64398
rect 2778 64152 2834 64161
rect 2778 64087 2834 64096
rect 2502 64016 2558 64025
rect 2502 63951 2504 63960
rect 2556 63951 2558 63960
rect 2780 63980 2832 63986
rect 2504 63922 2556 63928
rect 2884 63968 2912 64398
rect 2976 63986 3004 64466
rect 3068 64462 3096 67118
rect 3528 67046 3556 73170
rect 3608 72276 3660 72282
rect 3608 72218 3660 72224
rect 3516 67040 3568 67046
rect 3516 66982 3568 66988
rect 3516 66632 3568 66638
rect 3516 66574 3568 66580
rect 3240 65612 3292 65618
rect 3240 65554 3292 65560
rect 3056 64456 3108 64462
rect 3056 64398 3108 64404
rect 2832 63940 2912 63968
rect 2964 63980 3016 63986
rect 2780 63922 2832 63928
rect 2964 63922 3016 63928
rect 2582 63676 2890 63696
rect 2582 63674 2588 63676
rect 2644 63674 2668 63676
rect 2724 63674 2748 63676
rect 2804 63674 2828 63676
rect 2884 63674 2890 63676
rect 2644 63622 2646 63674
rect 2826 63622 2828 63674
rect 2582 63620 2588 63622
rect 2644 63620 2668 63622
rect 2724 63620 2748 63622
rect 2804 63620 2828 63622
rect 2884 63620 2890 63622
rect 2582 63600 2890 63620
rect 2504 63572 2556 63578
rect 2504 63514 2556 63520
rect 2412 62484 2464 62490
rect 2412 62426 2464 62432
rect 2332 62342 2452 62370
rect 2318 61976 2374 61985
rect 2318 61911 2374 61920
rect 2332 61810 2360 61911
rect 2320 61804 2372 61810
rect 2320 61746 2372 61752
rect 2320 61192 2372 61198
rect 2320 61134 2372 61140
rect 2226 59392 2282 59401
rect 2226 59327 2282 59336
rect 2148 59214 2268 59242
rect 2136 59152 2188 59158
rect 2136 59094 2188 59100
rect 2044 56772 2096 56778
rect 2044 56714 2096 56720
rect 1860 56704 1912 56710
rect 1860 56646 1912 56652
rect 1952 56704 2004 56710
rect 1952 56646 2004 56652
rect 1860 56160 1912 56166
rect 1860 56102 1912 56108
rect 1872 55282 1900 56102
rect 1860 55276 1912 55282
rect 1860 55218 1912 55224
rect 1964 54482 1992 56646
rect 2044 55276 2096 55282
rect 2044 55218 2096 55224
rect 1872 54454 1992 54482
rect 1768 49972 1820 49978
rect 1768 49914 1820 49920
rect 1768 49836 1820 49842
rect 1768 49778 1820 49784
rect 1490 49736 1546 49745
rect 1490 49671 1492 49680
rect 1544 49671 1546 49680
rect 1492 49642 1544 49648
rect 1490 49192 1546 49201
rect 1490 49127 1546 49136
rect 1504 49094 1532 49127
rect 1492 49088 1544 49094
rect 1492 49030 1544 49036
rect 1490 48648 1546 48657
rect 1490 48583 1492 48592
rect 1544 48583 1546 48592
rect 1492 48554 1544 48560
rect 1490 48104 1546 48113
rect 1490 48039 1546 48048
rect 1504 48006 1532 48039
rect 1492 48000 1544 48006
rect 1492 47942 1544 47948
rect 1676 47660 1728 47666
rect 1676 47602 1728 47608
rect 1490 47560 1546 47569
rect 1490 47495 1492 47504
rect 1544 47495 1546 47504
rect 1492 47466 1544 47472
rect 1492 47184 1544 47190
rect 1492 47126 1544 47132
rect 1504 47025 1532 47126
rect 1490 47016 1546 47025
rect 1490 46951 1546 46960
rect 1584 46572 1636 46578
rect 1584 46514 1636 46520
rect 1492 46368 1544 46374
rect 1490 46336 1492 46345
rect 1544 46336 1546 46345
rect 1490 46271 1546 46280
rect 1492 45824 1544 45830
rect 1490 45792 1492 45801
rect 1544 45792 1546 45801
rect 1490 45727 1546 45736
rect 1320 45526 1440 45554
rect 1320 41818 1348 45526
rect 1400 45484 1452 45490
rect 1400 45426 1452 45432
rect 1412 42362 1440 45426
rect 1492 45280 1544 45286
rect 1490 45248 1492 45257
rect 1544 45248 1546 45257
rect 1490 45183 1546 45192
rect 1492 44736 1544 44742
rect 1490 44704 1492 44713
rect 1544 44704 1546 44713
rect 1490 44639 1546 44648
rect 1492 44192 1544 44198
rect 1490 44160 1492 44169
rect 1544 44160 1546 44169
rect 1490 44095 1546 44104
rect 1492 43648 1544 43654
rect 1490 43616 1492 43625
rect 1544 43616 1546 43625
rect 1490 43551 1546 43560
rect 1492 43104 1544 43110
rect 1490 43072 1492 43081
rect 1544 43072 1546 43081
rect 1490 43007 1546 43016
rect 1492 42560 1544 42566
rect 1490 42528 1492 42537
rect 1544 42528 1546 42537
rect 1490 42463 1546 42472
rect 1400 42356 1452 42362
rect 1400 42298 1452 42304
rect 1400 42220 1452 42226
rect 1400 42162 1452 42168
rect 1308 41812 1360 41818
rect 1308 41754 1360 41760
rect 1308 41540 1360 41546
rect 1308 41482 1360 41488
rect 1320 41274 1348 41482
rect 1308 41268 1360 41274
rect 1308 41210 1360 41216
rect 1412 41120 1440 42162
rect 1492 42016 1544 42022
rect 1490 41984 1492 41993
rect 1544 41984 1546 41993
rect 1490 41919 1546 41928
rect 1492 41472 1544 41478
rect 1490 41440 1492 41449
rect 1544 41440 1546 41449
rect 1490 41375 1546 41384
rect 1492 41268 1544 41274
rect 1492 41210 1544 41216
rect 1320 41092 1440 41120
rect 1320 38894 1348 41092
rect 1504 41018 1532 41210
rect 1412 40990 1532 41018
rect 1412 40730 1440 40990
rect 1492 40928 1544 40934
rect 1490 40896 1492 40905
rect 1544 40896 1546 40905
rect 1490 40831 1546 40840
rect 1400 40724 1452 40730
rect 1400 40666 1452 40672
rect 1596 40610 1624 46514
rect 1412 40582 1624 40610
rect 1412 40202 1440 40582
rect 1584 40520 1636 40526
rect 1584 40462 1636 40468
rect 1492 40384 1544 40390
rect 1490 40352 1492 40361
rect 1544 40352 1546 40361
rect 1490 40287 1546 40296
rect 1412 40174 1532 40202
rect 1400 40044 1452 40050
rect 1400 39986 1452 39992
rect 1412 39681 1440 39986
rect 1398 39672 1454 39681
rect 1398 39607 1454 39616
rect 1400 39432 1452 39438
rect 1400 39374 1452 39380
rect 1412 39137 1440 39374
rect 1398 39128 1454 39137
rect 1398 39063 1454 39072
rect 1400 38956 1452 38962
rect 1400 38898 1452 38904
rect 1308 38888 1360 38894
rect 1308 38830 1360 38836
rect 1412 38593 1440 38898
rect 1398 38584 1454 38593
rect 1398 38519 1454 38528
rect 1308 38412 1360 38418
rect 1308 38354 1360 38360
rect 1320 37398 1348 38354
rect 1400 38344 1452 38350
rect 1400 38286 1452 38292
rect 1412 38049 1440 38286
rect 1398 38040 1454 38049
rect 1398 37975 1454 37984
rect 1400 37868 1452 37874
rect 1400 37810 1452 37816
rect 1412 37505 1440 37810
rect 1398 37496 1454 37505
rect 1398 37431 1454 37440
rect 1308 37392 1360 37398
rect 1308 37334 1360 37340
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 1412 36961 1440 37198
rect 1398 36952 1454 36961
rect 1398 36887 1454 36896
rect 1400 36780 1452 36786
rect 1400 36722 1452 36728
rect 1412 36417 1440 36722
rect 1398 36408 1454 36417
rect 1398 36343 1454 36352
rect 1504 36310 1532 40174
rect 1492 36304 1544 36310
rect 1492 36246 1544 36252
rect 1400 36168 1452 36174
rect 1596 36122 1624 40462
rect 1400 36110 1452 36116
rect 1412 35873 1440 36110
rect 1504 36094 1624 36122
rect 1398 35864 1454 35873
rect 1398 35799 1454 35808
rect 1400 35692 1452 35698
rect 1400 35634 1452 35640
rect 1412 35329 1440 35634
rect 1398 35320 1454 35329
rect 1216 35284 1268 35290
rect 1398 35255 1454 35264
rect 1216 35226 1268 35232
rect 1400 35080 1452 35086
rect 1400 35022 1452 35028
rect 1412 34785 1440 35022
rect 1398 34776 1454 34785
rect 1398 34711 1454 34720
rect 1400 34604 1452 34610
rect 1400 34546 1452 34552
rect 1412 34241 1440 34546
rect 1398 34232 1454 34241
rect 1398 34167 1454 34176
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1412 33697 1440 33934
rect 1398 33688 1454 33697
rect 1398 33623 1454 33632
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1412 33017 1440 33458
rect 1398 33008 1454 33017
rect 1398 32943 1454 32952
rect 1400 32904 1452 32910
rect 1400 32846 1452 32852
rect 1412 32473 1440 32846
rect 1398 32464 1454 32473
rect 1308 32428 1360 32434
rect 1398 32399 1454 32408
rect 1308 32370 1360 32376
rect 1320 31929 1348 32370
rect 1306 31920 1362 31929
rect 1306 31855 1362 31864
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 31385 1440 31758
rect 1398 31376 1454 31385
rect 1308 31340 1360 31346
rect 1398 31311 1454 31320
rect 1308 31282 1360 31288
rect 1320 30841 1348 31282
rect 1306 30832 1362 30841
rect 1504 30802 1532 36094
rect 1584 36032 1636 36038
rect 1584 35974 1636 35980
rect 1596 33658 1624 35974
rect 1688 35834 1716 47602
rect 1780 39098 1808 49778
rect 1872 49434 1900 54454
rect 1952 53100 2004 53106
rect 1952 53042 2004 53048
rect 1860 49428 1912 49434
rect 1860 49370 1912 49376
rect 1860 49224 1912 49230
rect 1860 49166 1912 49172
rect 1872 44742 1900 49166
rect 1964 44826 1992 53042
rect 2056 45082 2084 55218
rect 2148 52154 2176 59094
rect 2240 58070 2268 59214
rect 2228 58064 2280 58070
rect 2228 58006 2280 58012
rect 2228 57928 2280 57934
rect 2228 57870 2280 57876
rect 2240 56710 2268 57870
rect 2228 56704 2280 56710
rect 2228 56646 2280 56652
rect 2332 56522 2360 61134
rect 2424 56658 2452 62342
rect 2516 57032 2544 63514
rect 2872 63436 2924 63442
rect 2872 63378 2924 63384
rect 2780 63368 2832 63374
rect 2780 63310 2832 63316
rect 2596 63232 2648 63238
rect 2596 63174 2648 63180
rect 2688 63232 2740 63238
rect 2688 63174 2740 63180
rect 2608 62830 2636 63174
rect 2596 62824 2648 62830
rect 2596 62766 2648 62772
rect 2700 62762 2728 63174
rect 2792 62801 2820 63310
rect 2884 62898 2912 63378
rect 2976 63034 3004 63922
rect 2964 63028 3016 63034
rect 2964 62970 3016 62976
rect 2872 62892 2924 62898
rect 2872 62834 2924 62840
rect 2778 62792 2834 62801
rect 2688 62756 2740 62762
rect 2778 62727 2834 62736
rect 2688 62698 2740 62704
rect 2582 62588 2890 62608
rect 2582 62586 2588 62588
rect 2644 62586 2668 62588
rect 2724 62586 2748 62588
rect 2804 62586 2828 62588
rect 2884 62586 2890 62588
rect 2644 62534 2646 62586
rect 2826 62534 2828 62586
rect 2582 62532 2588 62534
rect 2644 62532 2668 62534
rect 2724 62532 2748 62534
rect 2804 62532 2828 62534
rect 2884 62532 2890 62534
rect 2582 62512 2890 62532
rect 3252 62354 3280 65554
rect 3528 65550 3556 66574
rect 3620 66314 3648 72218
rect 3712 70854 3740 73630
rect 3792 72616 3844 72622
rect 3792 72558 3844 72564
rect 3976 72616 4028 72622
rect 3976 72558 4028 72564
rect 3804 71602 3832 72558
rect 3884 72072 3936 72078
rect 3884 72014 3936 72020
rect 3792 71596 3844 71602
rect 3792 71538 3844 71544
rect 3700 70848 3752 70854
rect 3700 70790 3752 70796
rect 3804 66638 3832 71538
rect 3896 70990 3924 72014
rect 3988 71058 4016 72558
rect 4080 72078 4108 74054
rect 4213 74012 4521 74032
rect 4213 74010 4219 74012
rect 4275 74010 4299 74012
rect 4355 74010 4379 74012
rect 4435 74010 4459 74012
rect 4515 74010 4521 74012
rect 4275 73958 4277 74010
rect 4457 73958 4459 74010
rect 4213 73956 4219 73958
rect 4275 73956 4299 73958
rect 4355 73956 4379 73958
rect 4435 73956 4459 73958
rect 4515 73956 4521 73958
rect 4213 73936 4521 73956
rect 4712 73840 4764 73846
rect 4712 73782 4764 73788
rect 4528 73772 4580 73778
rect 4528 73714 4580 73720
rect 4540 73234 4568 73714
rect 4528 73228 4580 73234
rect 4528 73170 4580 73176
rect 4213 72924 4521 72944
rect 4213 72922 4219 72924
rect 4275 72922 4299 72924
rect 4355 72922 4379 72924
rect 4435 72922 4459 72924
rect 4515 72922 4521 72924
rect 4275 72870 4277 72922
rect 4457 72870 4459 72922
rect 4213 72868 4219 72870
rect 4275 72868 4299 72870
rect 4355 72868 4379 72870
rect 4435 72868 4459 72870
rect 4515 72868 4521 72870
rect 4213 72848 4521 72868
rect 4068 72072 4120 72078
rect 4068 72014 4120 72020
rect 4213 71836 4521 71856
rect 4213 71834 4219 71836
rect 4275 71834 4299 71836
rect 4355 71834 4379 71836
rect 4435 71834 4459 71836
rect 4515 71834 4521 71836
rect 4275 71782 4277 71834
rect 4457 71782 4459 71834
rect 4213 71780 4219 71782
rect 4275 71780 4299 71782
rect 4355 71780 4379 71782
rect 4435 71780 4459 71782
rect 4515 71780 4521 71782
rect 4213 71760 4521 71780
rect 4620 71732 4672 71738
rect 4620 71674 4672 71680
rect 3976 71052 4028 71058
rect 3976 70994 4028 71000
rect 3884 70984 3936 70990
rect 3884 70926 3936 70932
rect 3884 70848 3936 70854
rect 3884 70790 3936 70796
rect 3792 66632 3844 66638
rect 3896 66609 3924 70790
rect 3792 66574 3844 66580
rect 3882 66600 3938 66609
rect 3882 66535 3938 66544
rect 3988 66484 4016 70994
rect 4213 70748 4521 70768
rect 4213 70746 4219 70748
rect 4275 70746 4299 70748
rect 4355 70746 4379 70748
rect 4435 70746 4459 70748
rect 4515 70746 4521 70748
rect 4275 70694 4277 70746
rect 4457 70694 4459 70746
rect 4213 70692 4219 70694
rect 4275 70692 4299 70694
rect 4355 70692 4379 70694
rect 4435 70692 4459 70694
rect 4515 70692 4521 70694
rect 4213 70672 4521 70692
rect 4213 69660 4521 69680
rect 4213 69658 4219 69660
rect 4275 69658 4299 69660
rect 4355 69658 4379 69660
rect 4435 69658 4459 69660
rect 4515 69658 4521 69660
rect 4275 69606 4277 69658
rect 4457 69606 4459 69658
rect 4213 69604 4219 69606
rect 4275 69604 4299 69606
rect 4355 69604 4379 69606
rect 4435 69604 4459 69606
rect 4515 69604 4521 69606
rect 4213 69584 4521 69604
rect 4213 68572 4521 68592
rect 4213 68570 4219 68572
rect 4275 68570 4299 68572
rect 4355 68570 4379 68572
rect 4435 68570 4459 68572
rect 4515 68570 4521 68572
rect 4275 68518 4277 68570
rect 4457 68518 4459 68570
rect 4213 68516 4219 68518
rect 4275 68516 4299 68518
rect 4355 68516 4379 68518
rect 4435 68516 4459 68518
rect 4515 68516 4521 68518
rect 4213 68496 4521 68516
rect 4213 67484 4521 67504
rect 4213 67482 4219 67484
rect 4275 67482 4299 67484
rect 4355 67482 4379 67484
rect 4435 67482 4459 67484
rect 4515 67482 4521 67484
rect 4275 67430 4277 67482
rect 4457 67430 4459 67482
rect 4213 67428 4219 67430
rect 4275 67428 4299 67430
rect 4355 67428 4379 67430
rect 4435 67428 4459 67430
rect 4515 67428 4521 67430
rect 4213 67408 4521 67428
rect 4068 67040 4120 67046
rect 4068 66982 4120 66988
rect 3804 66456 4016 66484
rect 3620 66286 3740 66314
rect 3712 66230 3740 66286
rect 3700 66224 3752 66230
rect 3700 66166 3752 66172
rect 3608 66156 3660 66162
rect 3608 66098 3660 66104
rect 3620 65754 3648 66098
rect 3608 65748 3660 65754
rect 3608 65690 3660 65696
rect 3804 65686 3832 66456
rect 3882 66328 3938 66337
rect 3882 66263 3938 66272
rect 3792 65680 3844 65686
rect 3792 65622 3844 65628
rect 3516 65544 3568 65550
rect 3516 65486 3568 65492
rect 3528 63442 3556 65486
rect 3332 63436 3384 63442
rect 3332 63378 3384 63384
rect 3516 63436 3568 63442
rect 3516 63378 3568 63384
rect 3240 62348 3292 62354
rect 3240 62290 3292 62296
rect 2582 61500 2890 61520
rect 2582 61498 2588 61500
rect 2644 61498 2668 61500
rect 2724 61498 2748 61500
rect 2804 61498 2828 61500
rect 2884 61498 2890 61500
rect 2644 61446 2646 61498
rect 2826 61446 2828 61498
rect 2582 61444 2588 61446
rect 2644 61444 2668 61446
rect 2724 61444 2748 61446
rect 2804 61444 2828 61446
rect 2884 61444 2890 61446
rect 2582 61424 2890 61444
rect 3252 60734 3280 62290
rect 3068 60706 3280 60734
rect 2582 60412 2890 60432
rect 2582 60410 2588 60412
rect 2644 60410 2668 60412
rect 2724 60410 2748 60412
rect 2804 60410 2828 60412
rect 2884 60410 2890 60412
rect 2644 60358 2646 60410
rect 2826 60358 2828 60410
rect 2582 60356 2588 60358
rect 2644 60356 2668 60358
rect 2724 60356 2748 60358
rect 2804 60356 2828 60358
rect 2884 60356 2890 60358
rect 2582 60336 2890 60356
rect 2582 59324 2890 59344
rect 2582 59322 2588 59324
rect 2644 59322 2668 59324
rect 2724 59322 2748 59324
rect 2804 59322 2828 59324
rect 2884 59322 2890 59324
rect 2644 59270 2646 59322
rect 2826 59270 2828 59322
rect 2582 59268 2588 59270
rect 2644 59268 2668 59270
rect 2724 59268 2748 59270
rect 2804 59268 2828 59270
rect 2884 59268 2890 59270
rect 2582 59248 2890 59268
rect 2582 58236 2890 58256
rect 2582 58234 2588 58236
rect 2644 58234 2668 58236
rect 2724 58234 2748 58236
rect 2804 58234 2828 58236
rect 2884 58234 2890 58236
rect 2644 58182 2646 58234
rect 2826 58182 2828 58234
rect 2582 58180 2588 58182
rect 2644 58180 2668 58182
rect 2724 58180 2748 58182
rect 2804 58180 2828 58182
rect 2884 58180 2890 58182
rect 2582 58160 2890 58180
rect 2596 57928 2648 57934
rect 2596 57870 2648 57876
rect 2608 57458 2636 57870
rect 2780 57792 2832 57798
rect 2780 57734 2832 57740
rect 2792 57497 2820 57734
rect 2778 57488 2834 57497
rect 2596 57452 2648 57458
rect 2778 57423 2834 57432
rect 2596 57394 2648 57400
rect 2964 57248 3016 57254
rect 2964 57190 3016 57196
rect 2582 57148 2890 57168
rect 2582 57146 2588 57148
rect 2644 57146 2668 57148
rect 2724 57146 2748 57148
rect 2804 57146 2828 57148
rect 2884 57146 2890 57148
rect 2644 57094 2646 57146
rect 2826 57094 2828 57146
rect 2582 57092 2588 57094
rect 2644 57092 2668 57094
rect 2724 57092 2748 57094
rect 2804 57092 2828 57094
rect 2884 57092 2890 57094
rect 2582 57072 2890 57092
rect 2516 57004 2636 57032
rect 2424 56630 2544 56658
rect 2332 56494 2452 56522
rect 2320 55752 2372 55758
rect 2320 55694 2372 55700
rect 2228 53576 2280 53582
rect 2228 53518 2280 53524
rect 2136 52148 2188 52154
rect 2136 52090 2188 52096
rect 2136 52012 2188 52018
rect 2136 51954 2188 51960
rect 2148 51474 2176 51954
rect 2240 51814 2268 53518
rect 2228 51808 2280 51814
rect 2228 51750 2280 51756
rect 2136 51468 2188 51474
rect 2136 51410 2188 51416
rect 2240 51406 2268 51750
rect 2332 51649 2360 55694
rect 2424 52698 2452 56494
rect 2412 52692 2464 52698
rect 2412 52634 2464 52640
rect 2516 52193 2544 56630
rect 2608 56506 2636 57004
rect 2688 56840 2740 56846
rect 2688 56782 2740 56788
rect 2596 56500 2648 56506
rect 2596 56442 2648 56448
rect 2700 56370 2728 56782
rect 2872 56704 2924 56710
rect 2872 56646 2924 56652
rect 2688 56364 2740 56370
rect 2688 56306 2740 56312
rect 2884 56302 2912 56646
rect 2872 56296 2924 56302
rect 2872 56238 2924 56244
rect 2582 56060 2890 56080
rect 2582 56058 2588 56060
rect 2644 56058 2668 56060
rect 2724 56058 2748 56060
rect 2804 56058 2828 56060
rect 2884 56058 2890 56060
rect 2644 56006 2646 56058
rect 2826 56006 2828 56058
rect 2582 56004 2588 56006
rect 2644 56004 2668 56006
rect 2724 56004 2748 56006
rect 2804 56004 2828 56006
rect 2884 56004 2890 56006
rect 2582 55984 2890 56004
rect 2976 55865 3004 57190
rect 3068 56370 3096 60706
rect 3240 60648 3292 60654
rect 3240 60590 3292 60596
rect 3148 57520 3200 57526
rect 3148 57462 3200 57468
rect 3160 56778 3188 57462
rect 3252 57202 3280 60590
rect 3344 57526 3372 63378
rect 3792 62212 3844 62218
rect 3792 62154 3844 62160
rect 3700 61736 3752 61742
rect 3700 61678 3752 61684
rect 3424 60104 3476 60110
rect 3424 60046 3476 60052
rect 3332 57520 3384 57526
rect 3332 57462 3384 57468
rect 3252 57174 3372 57202
rect 3240 57044 3292 57050
rect 3240 56986 3292 56992
rect 3148 56772 3200 56778
rect 3148 56714 3200 56720
rect 3056 56364 3108 56370
rect 3056 56306 3108 56312
rect 3054 56264 3110 56273
rect 3054 56199 3056 56208
rect 3108 56199 3110 56208
rect 3056 56170 3108 56176
rect 2962 55856 3018 55865
rect 2962 55791 3018 55800
rect 3056 55684 3108 55690
rect 3056 55626 3108 55632
rect 2688 55412 2740 55418
rect 2688 55354 2740 55360
rect 2964 55412 3016 55418
rect 2964 55354 3016 55360
rect 2700 55146 2728 55354
rect 2688 55140 2740 55146
rect 2688 55082 2740 55088
rect 2582 54972 2890 54992
rect 2582 54970 2588 54972
rect 2644 54970 2668 54972
rect 2724 54970 2748 54972
rect 2804 54970 2828 54972
rect 2884 54970 2890 54972
rect 2644 54918 2646 54970
rect 2826 54918 2828 54970
rect 2582 54916 2588 54918
rect 2644 54916 2668 54918
rect 2724 54916 2748 54918
rect 2804 54916 2828 54918
rect 2884 54916 2890 54918
rect 2582 54896 2890 54916
rect 2976 54777 3004 55354
rect 2962 54768 3018 54777
rect 2962 54703 3018 54712
rect 2964 54120 3016 54126
rect 2964 54062 3016 54068
rect 2582 53884 2890 53904
rect 2582 53882 2588 53884
rect 2644 53882 2668 53884
rect 2724 53882 2748 53884
rect 2804 53882 2828 53884
rect 2884 53882 2890 53884
rect 2644 53830 2646 53882
rect 2826 53830 2828 53882
rect 2582 53828 2588 53830
rect 2644 53828 2668 53830
rect 2724 53828 2748 53830
rect 2804 53828 2828 53830
rect 2884 53828 2890 53830
rect 2582 53808 2890 53828
rect 2780 53100 2832 53106
rect 2780 53042 2832 53048
rect 2792 53009 2820 53042
rect 2778 53000 2834 53009
rect 2778 52935 2834 52944
rect 2582 52796 2890 52816
rect 2582 52794 2588 52796
rect 2644 52794 2668 52796
rect 2724 52794 2748 52796
rect 2804 52794 2828 52796
rect 2884 52794 2890 52796
rect 2644 52742 2646 52794
rect 2826 52742 2828 52794
rect 2582 52740 2588 52742
rect 2644 52740 2668 52742
rect 2724 52740 2748 52742
rect 2804 52740 2828 52742
rect 2884 52740 2890 52742
rect 2582 52720 2890 52740
rect 2502 52184 2558 52193
rect 2502 52119 2558 52128
rect 2504 52012 2556 52018
rect 2504 51954 2556 51960
rect 2318 51640 2374 51649
rect 2318 51575 2374 51584
rect 2412 51604 2464 51610
rect 2412 51546 2464 51552
rect 2424 51513 2452 51546
rect 2410 51504 2466 51513
rect 2320 51468 2372 51474
rect 2410 51439 2466 51448
rect 2320 51410 2372 51416
rect 2228 51400 2280 51406
rect 2228 51342 2280 51348
rect 2136 51264 2188 51270
rect 2136 51206 2188 51212
rect 2148 46714 2176 51206
rect 2226 51096 2282 51105
rect 2226 51031 2282 51040
rect 2136 46708 2188 46714
rect 2136 46650 2188 46656
rect 2136 46572 2188 46578
rect 2136 46514 2188 46520
rect 2148 45966 2176 46514
rect 2240 46170 2268 51031
rect 2332 50998 2360 51410
rect 2412 51400 2464 51406
rect 2412 51342 2464 51348
rect 2424 51066 2452 51342
rect 2412 51060 2464 51066
rect 2412 51002 2464 51008
rect 2320 50992 2372 50998
rect 2320 50934 2372 50940
rect 2332 50318 2360 50934
rect 2412 50924 2464 50930
rect 2412 50866 2464 50872
rect 2320 50312 2372 50318
rect 2320 50254 2372 50260
rect 2320 48136 2372 48142
rect 2320 48078 2372 48084
rect 2228 46164 2280 46170
rect 2228 46106 2280 46112
rect 2136 45960 2188 45966
rect 2136 45902 2188 45908
rect 2044 45076 2096 45082
rect 2044 45018 2096 45024
rect 2148 44878 2176 45902
rect 2228 45892 2280 45898
rect 2228 45834 2280 45840
rect 2136 44872 2188 44878
rect 1964 44798 2084 44826
rect 2136 44814 2188 44820
rect 1860 44736 1912 44742
rect 1860 44678 1912 44684
rect 2056 44418 2084 44798
rect 2136 44736 2188 44742
rect 2136 44678 2188 44684
rect 1964 44390 2084 44418
rect 1860 42696 1912 42702
rect 1860 42638 1912 42644
rect 1768 39092 1820 39098
rect 1768 39034 1820 39040
rect 1768 38888 1820 38894
rect 1768 38830 1820 38836
rect 1676 35828 1728 35834
rect 1676 35770 1728 35776
rect 1780 35714 1808 38830
rect 1688 35686 1808 35714
rect 1584 33652 1636 33658
rect 1584 33594 1636 33600
rect 1688 33538 1716 35686
rect 1768 35012 1820 35018
rect 1768 34954 1820 34960
rect 1596 33510 1716 33538
rect 1306 30767 1362 30776
rect 1492 30796 1544 30802
rect 1492 30738 1544 30744
rect 1400 30728 1452 30734
rect 1596 30682 1624 33510
rect 1676 32292 1728 32298
rect 1676 32234 1728 32240
rect 1688 31482 1716 32234
rect 1676 31476 1728 31482
rect 1676 31418 1728 31424
rect 1676 31204 1728 31210
rect 1676 31146 1728 31152
rect 1400 30670 1452 30676
rect 1412 30297 1440 30670
rect 1504 30654 1624 30682
rect 1398 30288 1454 30297
rect 1308 30252 1360 30258
rect 1398 30223 1454 30232
rect 1308 30194 1360 30200
rect 1320 29753 1348 30194
rect 1306 29744 1362 29753
rect 1306 29679 1362 29688
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1412 29209 1440 29582
rect 1398 29200 1454 29209
rect 1308 29164 1360 29170
rect 1398 29135 1454 29144
rect 1308 29106 1360 29112
rect 1216 29096 1268 29102
rect 1216 29038 1268 29044
rect 1228 28150 1256 29038
rect 1320 28665 1348 29106
rect 1504 29050 1532 30654
rect 1584 30388 1636 30394
rect 1584 30330 1636 30336
rect 1596 29850 1624 30330
rect 1688 30122 1716 31146
rect 1780 30938 1808 34954
rect 1768 30932 1820 30938
rect 1768 30874 1820 30880
rect 1676 30116 1728 30122
rect 1676 30058 1728 30064
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 1768 29844 1820 29850
rect 1768 29786 1820 29792
rect 1676 29504 1728 29510
rect 1676 29446 1728 29452
rect 1688 29306 1716 29446
rect 1676 29300 1728 29306
rect 1676 29242 1728 29248
rect 1504 29022 1624 29050
rect 1492 28960 1544 28966
rect 1492 28902 1544 28908
rect 1306 28656 1362 28665
rect 1306 28591 1362 28600
rect 1400 28552 1452 28558
rect 1400 28494 1452 28500
rect 1216 28144 1268 28150
rect 1412 28121 1440 28494
rect 1216 28086 1268 28092
rect 1398 28112 1454 28121
rect 1308 28076 1360 28082
rect 1398 28047 1454 28056
rect 1308 28018 1360 28024
rect 1216 28008 1268 28014
rect 1216 27950 1268 27956
rect 1228 27146 1256 27950
rect 1320 27577 1348 28018
rect 1306 27568 1362 27577
rect 1306 27503 1362 27512
rect 1228 27118 1348 27146
rect 1216 27056 1268 27062
rect 1216 26998 1268 27004
rect 1124 12776 1176 12782
rect 1124 12718 1176 12724
rect 1228 11914 1256 26998
rect 1136 11886 1256 11914
rect 1136 6186 1164 11886
rect 1320 11778 1348 27118
rect 1504 21622 1532 28902
rect 1596 27946 1624 29022
rect 1780 28218 1808 29786
rect 1872 29306 1900 42638
rect 1964 41274 1992 44390
rect 2044 44328 2096 44334
rect 2044 44270 2096 44276
rect 1952 41268 2004 41274
rect 1952 41210 2004 41216
rect 1950 41168 2006 41177
rect 1950 41103 2006 41112
rect 1964 36922 1992 41103
rect 1952 36916 2004 36922
rect 1952 36858 2004 36864
rect 2056 31482 2084 44270
rect 2148 41721 2176 44678
rect 2134 41712 2190 41721
rect 2134 41647 2190 41656
rect 2136 41608 2188 41614
rect 2136 41550 2188 41556
rect 2148 41138 2176 41550
rect 2136 41132 2188 41138
rect 2136 41074 2188 41080
rect 2148 40526 2176 41074
rect 2136 40520 2188 40526
rect 2136 40462 2188 40468
rect 2136 39432 2188 39438
rect 2136 39374 2188 39380
rect 2148 38962 2176 39374
rect 2136 38956 2188 38962
rect 2136 38898 2188 38904
rect 2148 38350 2176 38898
rect 2136 38344 2188 38350
rect 2136 38286 2188 38292
rect 2136 36780 2188 36786
rect 2136 36722 2188 36728
rect 2148 36174 2176 36722
rect 2136 36168 2188 36174
rect 2136 36110 2188 36116
rect 2148 35698 2176 36110
rect 2136 35692 2188 35698
rect 2136 35634 2188 35640
rect 2240 32570 2268 45834
rect 2332 41313 2360 48078
rect 2318 41304 2374 41313
rect 2318 41239 2374 41248
rect 2318 41168 2374 41177
rect 2318 41103 2374 41112
rect 2332 38554 2360 41103
rect 2424 39642 2452 50866
rect 2516 50368 2544 51954
rect 2778 51912 2834 51921
rect 2778 51847 2780 51856
rect 2832 51847 2834 51856
rect 2780 51818 2832 51824
rect 2582 51708 2890 51728
rect 2582 51706 2588 51708
rect 2644 51706 2668 51708
rect 2724 51706 2748 51708
rect 2804 51706 2828 51708
rect 2884 51706 2890 51708
rect 2644 51654 2646 51706
rect 2826 51654 2828 51706
rect 2582 51652 2588 51654
rect 2644 51652 2668 51654
rect 2724 51652 2748 51654
rect 2804 51652 2828 51654
rect 2884 51652 2890 51654
rect 2582 51632 2890 51652
rect 2596 51536 2648 51542
rect 2596 51478 2648 51484
rect 2608 51377 2636 51478
rect 2976 51406 3004 54062
rect 3068 53650 3096 55626
rect 3160 54262 3188 56714
rect 3148 54256 3200 54262
rect 3148 54198 3200 54204
rect 3252 54194 3280 56986
rect 3240 54188 3292 54194
rect 3240 54130 3292 54136
rect 3148 54120 3200 54126
rect 3344 54074 3372 57174
rect 3148 54062 3200 54068
rect 3056 53644 3108 53650
rect 3056 53586 3108 53592
rect 3056 53440 3108 53446
rect 3056 53382 3108 53388
rect 3068 53106 3096 53382
rect 3056 53100 3108 53106
rect 3056 53042 3108 53048
rect 3160 52986 3188 54062
rect 3252 54046 3372 54074
rect 3252 53145 3280 54046
rect 3238 53136 3294 53145
rect 3238 53071 3294 53080
rect 3068 52958 3188 52986
rect 2964 51400 3016 51406
rect 2594 51368 2650 51377
rect 2964 51342 3016 51348
rect 2594 51303 2650 51312
rect 3068 51074 3096 52958
rect 3240 52896 3292 52902
rect 3146 52864 3202 52873
rect 3240 52838 3292 52844
rect 3146 52799 3202 52808
rect 3160 52562 3188 52799
rect 3148 52556 3200 52562
rect 3148 52498 3200 52504
rect 3252 52494 3280 52838
rect 3240 52488 3292 52494
rect 3240 52430 3292 52436
rect 3148 52352 3200 52358
rect 3148 52294 3200 52300
rect 2976 51046 3096 51074
rect 2778 50824 2834 50833
rect 2778 50759 2780 50768
rect 2832 50759 2834 50768
rect 2780 50730 2832 50736
rect 2582 50620 2890 50640
rect 2582 50618 2588 50620
rect 2644 50618 2668 50620
rect 2724 50618 2748 50620
rect 2804 50618 2828 50620
rect 2884 50618 2890 50620
rect 2644 50566 2646 50618
rect 2826 50566 2828 50618
rect 2582 50564 2588 50566
rect 2644 50564 2668 50566
rect 2724 50564 2748 50566
rect 2804 50564 2828 50566
rect 2884 50564 2890 50566
rect 2582 50544 2890 50564
rect 2516 50340 2636 50368
rect 2502 50280 2558 50289
rect 2502 50215 2558 50224
rect 2516 50182 2544 50215
rect 2504 50176 2556 50182
rect 2504 50118 2556 50124
rect 2608 49688 2636 50340
rect 2516 49660 2636 49688
rect 2516 45558 2544 49660
rect 2582 49532 2890 49552
rect 2582 49530 2588 49532
rect 2644 49530 2668 49532
rect 2724 49530 2748 49532
rect 2804 49530 2828 49532
rect 2884 49530 2890 49532
rect 2644 49478 2646 49530
rect 2826 49478 2828 49530
rect 2582 49476 2588 49478
rect 2644 49476 2668 49478
rect 2724 49476 2748 49478
rect 2804 49476 2828 49478
rect 2884 49476 2890 49478
rect 2582 49456 2890 49476
rect 2582 48444 2890 48464
rect 2582 48442 2588 48444
rect 2644 48442 2668 48444
rect 2724 48442 2748 48444
rect 2804 48442 2828 48444
rect 2884 48442 2890 48444
rect 2644 48390 2646 48442
rect 2826 48390 2828 48442
rect 2582 48388 2588 48390
rect 2644 48388 2668 48390
rect 2724 48388 2748 48390
rect 2804 48388 2828 48390
rect 2884 48388 2890 48390
rect 2582 48368 2890 48388
rect 2582 47356 2890 47376
rect 2582 47354 2588 47356
rect 2644 47354 2668 47356
rect 2724 47354 2748 47356
rect 2804 47354 2828 47356
rect 2884 47354 2890 47356
rect 2644 47302 2646 47354
rect 2826 47302 2828 47354
rect 2582 47300 2588 47302
rect 2644 47300 2668 47302
rect 2724 47300 2748 47302
rect 2804 47300 2828 47302
rect 2884 47300 2890 47302
rect 2582 47280 2890 47300
rect 2582 46268 2890 46288
rect 2582 46266 2588 46268
rect 2644 46266 2668 46268
rect 2724 46266 2748 46268
rect 2804 46266 2828 46268
rect 2884 46266 2890 46268
rect 2644 46214 2646 46266
rect 2826 46214 2828 46266
rect 2582 46212 2588 46214
rect 2644 46212 2668 46214
rect 2724 46212 2748 46214
rect 2804 46212 2828 46214
rect 2884 46212 2890 46214
rect 2582 46192 2890 46212
rect 2686 46064 2742 46073
rect 2686 45999 2742 46008
rect 2596 45892 2648 45898
rect 2596 45834 2648 45840
rect 2504 45552 2556 45558
rect 2504 45494 2556 45500
rect 2608 45490 2636 45834
rect 2596 45484 2648 45490
rect 2596 45426 2648 45432
rect 2608 45336 2636 45426
rect 2700 45422 2728 45999
rect 2688 45416 2740 45422
rect 2688 45358 2740 45364
rect 2516 45308 2636 45336
rect 2516 44946 2544 45308
rect 2582 45180 2890 45200
rect 2582 45178 2588 45180
rect 2644 45178 2668 45180
rect 2724 45178 2748 45180
rect 2804 45178 2828 45180
rect 2884 45178 2890 45180
rect 2644 45126 2646 45178
rect 2826 45126 2828 45178
rect 2582 45124 2588 45126
rect 2644 45124 2668 45126
rect 2724 45124 2748 45126
rect 2804 45124 2828 45126
rect 2884 45124 2890 45126
rect 2582 45104 2890 45124
rect 2976 45082 3004 51046
rect 3056 50856 3108 50862
rect 3056 50798 3108 50804
rect 3068 50522 3096 50798
rect 3056 50516 3108 50522
rect 3056 50458 3108 50464
rect 3056 50312 3108 50318
rect 3056 50254 3108 50260
rect 3068 45966 3096 50254
rect 3056 45960 3108 45966
rect 3056 45902 3108 45908
rect 3160 45506 3188 52294
rect 3238 52184 3294 52193
rect 3436 52154 3464 60046
rect 3608 59628 3660 59634
rect 3608 59570 3660 59576
rect 3516 57452 3568 57458
rect 3516 57394 3568 57400
rect 3528 54126 3556 57394
rect 3620 56506 3648 59570
rect 3608 56500 3660 56506
rect 3608 56442 3660 56448
rect 3608 56364 3660 56370
rect 3608 56306 3660 56312
rect 3516 54120 3568 54126
rect 3516 54062 3568 54068
rect 3516 53032 3568 53038
rect 3516 52974 3568 52980
rect 3528 52442 3556 52974
rect 3620 52578 3648 56306
rect 3712 52698 3740 61678
rect 3804 53242 3832 62154
rect 3896 57050 3924 66263
rect 3976 66156 4028 66162
rect 3976 66098 4028 66104
rect 3988 65618 4016 66098
rect 3976 65612 4028 65618
rect 3976 65554 4028 65560
rect 3976 63368 4028 63374
rect 3976 63310 4028 63316
rect 3988 63073 4016 63310
rect 3974 63064 4030 63073
rect 3974 62999 4030 63008
rect 3884 57044 3936 57050
rect 3884 56986 3936 56992
rect 3884 56840 3936 56846
rect 3884 56782 3936 56788
rect 3792 53236 3844 53242
rect 3792 53178 3844 53184
rect 3700 52692 3752 52698
rect 3700 52634 3752 52640
rect 3620 52550 3832 52578
rect 3528 52414 3740 52442
rect 3608 52352 3660 52358
rect 3514 52320 3570 52329
rect 3608 52294 3660 52300
rect 3514 52255 3570 52264
rect 3238 52119 3294 52128
rect 3424 52148 3476 52154
rect 3252 51406 3280 52119
rect 3424 52090 3476 52096
rect 3424 51944 3476 51950
rect 3424 51886 3476 51892
rect 3240 51400 3292 51406
rect 3240 51342 3292 51348
rect 3240 51264 3292 51270
rect 3240 51206 3292 51212
rect 3252 45529 3280 51206
rect 3436 51074 3464 51886
rect 3344 51046 3464 51074
rect 3344 50794 3372 51046
rect 3528 50912 3556 52255
rect 3620 51066 3648 52294
rect 3608 51060 3660 51066
rect 3608 51002 3660 51008
rect 3436 50884 3556 50912
rect 3332 50788 3384 50794
rect 3332 50730 3384 50736
rect 3344 49706 3372 50730
rect 3436 50386 3464 50884
rect 3514 50824 3570 50833
rect 3514 50759 3570 50768
rect 3424 50380 3476 50386
rect 3424 50322 3476 50328
rect 3424 50244 3476 50250
rect 3424 50186 3476 50192
rect 3332 49700 3384 49706
rect 3332 49642 3384 49648
rect 3344 49162 3372 49642
rect 3332 49156 3384 49162
rect 3332 49098 3384 49104
rect 3344 47666 3372 49098
rect 3332 47660 3384 47666
rect 3332 47602 3384 47608
rect 3332 47048 3384 47054
rect 3332 46990 3384 46996
rect 3068 45478 3188 45506
rect 3238 45520 3294 45529
rect 2964 45076 3016 45082
rect 2964 45018 3016 45024
rect 2504 44940 2556 44946
rect 2504 44882 2556 44888
rect 2780 44736 2832 44742
rect 2780 44678 2832 44684
rect 2792 44282 2820 44678
rect 2792 44254 3004 44282
rect 2582 44092 2890 44112
rect 2582 44090 2588 44092
rect 2644 44090 2668 44092
rect 2724 44090 2748 44092
rect 2804 44090 2828 44092
rect 2884 44090 2890 44092
rect 2644 44038 2646 44090
rect 2826 44038 2828 44090
rect 2582 44036 2588 44038
rect 2644 44036 2668 44038
rect 2724 44036 2748 44038
rect 2804 44036 2828 44038
rect 2884 44036 2890 44038
rect 2582 44016 2890 44036
rect 2504 43784 2556 43790
rect 2504 43726 2556 43732
rect 2516 41698 2544 43726
rect 2582 43004 2890 43024
rect 2582 43002 2588 43004
rect 2644 43002 2668 43004
rect 2724 43002 2748 43004
rect 2804 43002 2828 43004
rect 2884 43002 2890 43004
rect 2644 42950 2646 43002
rect 2826 42950 2828 43002
rect 2582 42948 2588 42950
rect 2644 42948 2668 42950
rect 2724 42948 2748 42950
rect 2804 42948 2828 42950
rect 2884 42948 2890 42950
rect 2582 42928 2890 42948
rect 2582 41916 2890 41936
rect 2582 41914 2588 41916
rect 2644 41914 2668 41916
rect 2724 41914 2748 41916
rect 2804 41914 2828 41916
rect 2884 41914 2890 41916
rect 2644 41862 2646 41914
rect 2826 41862 2828 41914
rect 2582 41860 2588 41862
rect 2644 41860 2668 41862
rect 2724 41860 2748 41862
rect 2804 41860 2828 41862
rect 2884 41860 2890 41862
rect 2582 41840 2890 41860
rect 2516 41670 2636 41698
rect 2502 41576 2558 41585
rect 2502 41511 2558 41520
rect 2516 41177 2544 41511
rect 2502 41168 2558 41177
rect 2502 41103 2558 41112
rect 2608 41018 2636 41670
rect 2780 41608 2832 41614
rect 2780 41550 2832 41556
rect 2688 41540 2740 41546
rect 2688 41482 2740 41488
rect 2700 41138 2728 41482
rect 2792 41177 2820 41550
rect 2778 41168 2834 41177
rect 2688 41132 2740 41138
rect 2778 41103 2834 41112
rect 2688 41074 2740 41080
rect 2516 40990 2636 41018
rect 2412 39636 2464 39642
rect 2412 39578 2464 39584
rect 2412 39500 2464 39506
rect 2412 39442 2464 39448
rect 2320 38548 2372 38554
rect 2320 38490 2372 38496
rect 2320 37800 2372 37806
rect 2320 37742 2372 37748
rect 2332 37330 2360 37742
rect 2320 37324 2372 37330
rect 2320 37266 2372 37272
rect 2228 32564 2280 32570
rect 2228 32506 2280 32512
rect 2136 32428 2188 32434
rect 2136 32370 2188 32376
rect 2148 31822 2176 32370
rect 2424 32026 2452 39442
rect 2412 32020 2464 32026
rect 2412 31962 2464 31968
rect 2136 31816 2188 31822
rect 2136 31758 2188 31764
rect 2044 31476 2096 31482
rect 2044 31418 2096 31424
rect 2148 31346 2176 31758
rect 2516 31754 2544 40990
rect 2582 40828 2890 40848
rect 2582 40826 2588 40828
rect 2644 40826 2668 40828
rect 2724 40826 2748 40828
rect 2804 40826 2828 40828
rect 2884 40826 2890 40828
rect 2644 40774 2646 40826
rect 2826 40774 2828 40826
rect 2582 40772 2588 40774
rect 2644 40772 2668 40774
rect 2724 40772 2748 40774
rect 2804 40772 2828 40774
rect 2884 40772 2890 40774
rect 2582 40752 2890 40772
rect 2872 40520 2924 40526
rect 2872 40462 2924 40468
rect 2594 40080 2650 40089
rect 2884 40050 2912 40462
rect 2594 40015 2596 40024
rect 2648 40015 2650 40024
rect 2872 40044 2924 40050
rect 2596 39986 2648 39992
rect 2872 39986 2924 39992
rect 2582 39740 2890 39760
rect 2582 39738 2588 39740
rect 2644 39738 2668 39740
rect 2724 39738 2748 39740
rect 2804 39738 2828 39740
rect 2884 39738 2890 39740
rect 2644 39686 2646 39738
rect 2826 39686 2828 39738
rect 2582 39684 2588 39686
rect 2644 39684 2668 39686
rect 2724 39684 2748 39686
rect 2804 39684 2828 39686
rect 2884 39684 2890 39686
rect 2582 39664 2890 39684
rect 2582 38652 2890 38672
rect 2582 38650 2588 38652
rect 2644 38650 2668 38652
rect 2724 38650 2748 38652
rect 2804 38650 2828 38652
rect 2884 38650 2890 38652
rect 2644 38598 2646 38650
rect 2826 38598 2828 38650
rect 2582 38596 2588 38598
rect 2644 38596 2668 38598
rect 2724 38596 2748 38598
rect 2804 38596 2828 38598
rect 2884 38596 2890 38598
rect 2582 38576 2890 38596
rect 2780 38344 2832 38350
rect 2780 38286 2832 38292
rect 2792 37874 2820 38286
rect 2780 37868 2832 37874
rect 2780 37810 2832 37816
rect 2582 37564 2890 37584
rect 2582 37562 2588 37564
rect 2644 37562 2668 37564
rect 2724 37562 2748 37564
rect 2804 37562 2828 37564
rect 2884 37562 2890 37564
rect 2644 37510 2646 37562
rect 2826 37510 2828 37562
rect 2582 37508 2588 37510
rect 2644 37508 2668 37510
rect 2724 37508 2748 37510
rect 2804 37508 2828 37510
rect 2884 37508 2890 37510
rect 2582 37488 2890 37508
rect 2688 37256 2740 37262
rect 2688 37198 2740 37204
rect 2700 36854 2728 37198
rect 2688 36848 2740 36854
rect 2688 36790 2740 36796
rect 2582 36476 2890 36496
rect 2582 36474 2588 36476
rect 2644 36474 2668 36476
rect 2724 36474 2748 36476
rect 2804 36474 2828 36476
rect 2884 36474 2890 36476
rect 2644 36422 2646 36474
rect 2826 36422 2828 36474
rect 2582 36420 2588 36422
rect 2644 36420 2668 36422
rect 2724 36420 2748 36422
rect 2804 36420 2828 36422
rect 2884 36420 2890 36422
rect 2582 36400 2890 36420
rect 2582 35388 2890 35408
rect 2582 35386 2588 35388
rect 2644 35386 2668 35388
rect 2724 35386 2748 35388
rect 2804 35386 2828 35388
rect 2884 35386 2890 35388
rect 2644 35334 2646 35386
rect 2826 35334 2828 35386
rect 2582 35332 2588 35334
rect 2644 35332 2668 35334
rect 2724 35332 2748 35334
rect 2804 35332 2828 35334
rect 2884 35332 2890 35334
rect 2582 35312 2890 35332
rect 2582 34300 2890 34320
rect 2582 34298 2588 34300
rect 2644 34298 2668 34300
rect 2724 34298 2748 34300
rect 2804 34298 2828 34300
rect 2884 34298 2890 34300
rect 2644 34246 2646 34298
rect 2826 34246 2828 34298
rect 2582 34244 2588 34246
rect 2644 34244 2668 34246
rect 2724 34244 2748 34246
rect 2804 34244 2828 34246
rect 2884 34244 2890 34246
rect 2582 34224 2890 34244
rect 2582 33212 2890 33232
rect 2582 33210 2588 33212
rect 2644 33210 2668 33212
rect 2724 33210 2748 33212
rect 2804 33210 2828 33212
rect 2884 33210 2890 33212
rect 2644 33158 2646 33210
rect 2826 33158 2828 33210
rect 2582 33156 2588 33158
rect 2644 33156 2668 33158
rect 2724 33156 2748 33158
rect 2804 33156 2828 33158
rect 2884 33156 2890 33158
rect 2582 33136 2890 33156
rect 2582 32124 2890 32144
rect 2582 32122 2588 32124
rect 2644 32122 2668 32124
rect 2724 32122 2748 32124
rect 2804 32122 2828 32124
rect 2884 32122 2890 32124
rect 2644 32070 2646 32122
rect 2826 32070 2828 32122
rect 2582 32068 2588 32070
rect 2644 32068 2668 32070
rect 2724 32068 2748 32070
rect 2804 32068 2828 32070
rect 2884 32068 2890 32070
rect 2582 32048 2890 32068
rect 2424 31726 2544 31754
rect 2136 31340 2188 31346
rect 2136 31282 2188 31288
rect 1952 30796 2004 30802
rect 1952 30738 2004 30744
rect 1860 29300 1912 29306
rect 1860 29242 1912 29248
rect 1964 28762 1992 30738
rect 2148 30734 2176 31282
rect 2424 30938 2452 31726
rect 2582 31036 2890 31056
rect 2582 31034 2588 31036
rect 2644 31034 2668 31036
rect 2724 31034 2748 31036
rect 2804 31034 2828 31036
rect 2884 31034 2890 31036
rect 2644 30982 2646 31034
rect 2826 30982 2828 31034
rect 2582 30980 2588 30982
rect 2644 30980 2668 30982
rect 2724 30980 2748 30982
rect 2804 30980 2828 30982
rect 2884 30980 2890 30982
rect 2582 30960 2890 30980
rect 2976 30938 3004 44254
rect 3068 41154 3096 45478
rect 3238 45455 3294 45464
rect 3344 45336 3372 46990
rect 3160 45308 3372 45336
rect 3160 41274 3188 45308
rect 3238 45112 3294 45121
rect 3238 45047 3294 45056
rect 3148 41268 3200 41274
rect 3148 41210 3200 41216
rect 3068 41126 3188 41154
rect 3054 40080 3110 40089
rect 3054 40015 3110 40024
rect 3068 37806 3096 40015
rect 3160 39098 3188 41126
rect 3148 39092 3200 39098
rect 3148 39034 3200 39040
rect 3056 37800 3108 37806
rect 3056 37742 3108 37748
rect 3056 37188 3108 37194
rect 3056 37130 3108 37136
rect 2412 30932 2464 30938
rect 2412 30874 2464 30880
rect 2964 30932 3016 30938
rect 2964 30874 3016 30880
rect 2136 30728 2188 30734
rect 2136 30670 2188 30676
rect 2504 30728 2556 30734
rect 2504 30670 2556 30676
rect 2320 30252 2372 30258
rect 2320 30194 2372 30200
rect 2332 29714 2360 30194
rect 2516 29714 2544 30670
rect 2964 30184 3016 30190
rect 2964 30126 3016 30132
rect 2582 29948 2890 29968
rect 2582 29946 2588 29948
rect 2644 29946 2668 29948
rect 2724 29946 2748 29948
rect 2804 29946 2828 29948
rect 2884 29946 2890 29948
rect 2644 29894 2646 29946
rect 2826 29894 2828 29946
rect 2582 29892 2588 29894
rect 2644 29892 2668 29894
rect 2724 29892 2748 29894
rect 2804 29892 2828 29894
rect 2884 29892 2890 29894
rect 2582 29872 2890 29892
rect 2320 29708 2372 29714
rect 2320 29650 2372 29656
rect 2504 29708 2556 29714
rect 2504 29650 2556 29656
rect 2976 29238 3004 30126
rect 2964 29232 3016 29238
rect 2964 29174 3016 29180
rect 2044 28960 2096 28966
rect 2044 28902 2096 28908
rect 1952 28756 2004 28762
rect 1952 28698 2004 28704
rect 1768 28212 1820 28218
rect 1768 28154 1820 28160
rect 1584 27940 1636 27946
rect 1584 27882 1636 27888
rect 2056 27690 2084 28902
rect 2582 28860 2890 28880
rect 2582 28858 2588 28860
rect 2644 28858 2668 28860
rect 2724 28858 2748 28860
rect 2804 28858 2828 28860
rect 2884 28858 2890 28860
rect 2644 28806 2646 28858
rect 2826 28806 2828 28858
rect 2582 28804 2588 28806
rect 2644 28804 2668 28806
rect 2724 28804 2748 28806
rect 2804 28804 2828 28806
rect 2884 28804 2890 28806
rect 2582 28784 2890 28804
rect 2976 28642 3004 29174
rect 2884 28614 3004 28642
rect 2884 28558 2912 28614
rect 2872 28552 2924 28558
rect 2872 28494 2924 28500
rect 2504 28416 2556 28422
rect 2504 28358 2556 28364
rect 1964 27662 2084 27690
rect 2516 27674 2544 28358
rect 2884 28082 2912 28494
rect 2872 28076 2924 28082
rect 2872 28018 2924 28024
rect 2582 27772 2890 27792
rect 2582 27770 2588 27772
rect 2644 27770 2668 27772
rect 2724 27770 2748 27772
rect 2804 27770 2828 27772
rect 2884 27770 2890 27772
rect 2644 27718 2646 27770
rect 2826 27718 2828 27770
rect 2582 27716 2588 27718
rect 2644 27716 2668 27718
rect 2724 27716 2748 27718
rect 2804 27716 2828 27718
rect 2884 27716 2890 27718
rect 2582 27696 2890 27716
rect 2504 27668 2556 27674
rect 1964 27554 1992 27662
rect 2504 27610 2556 27616
rect 1872 27526 1992 27554
rect 2044 27600 2096 27606
rect 2044 27542 2096 27548
rect 1872 24410 1900 27526
rect 1952 27396 2004 27402
rect 1952 27338 2004 27344
rect 1964 27033 1992 27338
rect 1950 27024 2006 27033
rect 1950 26959 2006 26968
rect 1950 26344 2006 26353
rect 1950 26279 1952 26288
rect 2004 26279 2006 26288
rect 1952 26250 2004 26256
rect 1952 25900 2004 25906
rect 1952 25842 2004 25848
rect 1964 25809 1992 25842
rect 1950 25800 2006 25809
rect 1950 25735 2006 25744
rect 1950 25256 2006 25265
rect 1950 25191 1952 25200
rect 2004 25191 2006 25200
rect 1952 25162 2004 25168
rect 1952 24812 2004 24818
rect 1952 24754 2004 24760
rect 1964 24721 1992 24754
rect 1950 24712 2006 24721
rect 1950 24647 2006 24656
rect 1860 24404 1912 24410
rect 1860 24346 1912 24352
rect 1950 24168 2006 24177
rect 1950 24103 1952 24112
rect 2004 24103 2006 24112
rect 1952 24074 2004 24080
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1492 21616 1544 21622
rect 1492 21558 1544 21564
rect 1490 21448 1546 21457
rect 1490 21383 1492 21392
rect 1544 21383 1546 21392
rect 1492 21354 1544 21360
rect 1490 20904 1546 20913
rect 1490 20839 1546 20848
rect 1504 20806 1532 20839
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1490 20360 1546 20369
rect 1490 20295 1492 20304
rect 1544 20295 1546 20304
rect 1492 20266 1544 20272
rect 1688 19854 1716 22918
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1492 19712 1544 19718
rect 1490 19680 1492 19689
rect 1544 19680 1546 19689
rect 1490 19615 1546 19624
rect 1492 19168 1544 19174
rect 1490 19136 1492 19145
rect 1544 19136 1546 19145
rect 1490 19071 1546 19080
rect 1780 18766 1808 24006
rect 2056 23798 2084 27542
rect 2504 27532 2556 27538
rect 2504 27474 2556 27480
rect 2320 27464 2372 27470
rect 2320 27406 2372 27412
rect 2044 23792 2096 23798
rect 2044 23734 2096 23740
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 23633 1900 23666
rect 1858 23624 1914 23633
rect 1858 23559 1914 23568
rect 1950 23080 2006 23089
rect 1950 23015 1952 23024
rect 2004 23015 2006 23024
rect 1952 22986 2004 22992
rect 1952 22636 2004 22642
rect 1952 22578 2004 22584
rect 1964 22545 1992 22578
rect 1950 22536 2006 22545
rect 1950 22471 2006 22480
rect 1952 22024 2004 22030
rect 1950 21992 1952 22001
rect 2004 21992 2006 22001
rect 1950 21927 2006 21936
rect 1952 21888 2004 21894
rect 1952 21830 2004 21836
rect 1964 20466 1992 21830
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 2044 19440 2096 19446
rect 2044 19382 2096 19388
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1492 18624 1544 18630
rect 1490 18592 1492 18601
rect 1544 18592 1546 18601
rect 1490 18527 1546 18536
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1676 18080 1728 18086
rect 1544 18048 1546 18057
rect 1676 18022 1728 18028
rect 1490 17983 1546 17992
rect 1492 17536 1544 17542
rect 1490 17504 1492 17513
rect 1544 17504 1546 17513
rect 1490 17439 1546 17448
rect 1688 17202 1716 18022
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1492 16992 1544 16998
rect 1490 16960 1492 16969
rect 1676 16992 1728 16998
rect 1544 16960 1546 16969
rect 1676 16934 1728 16940
rect 1490 16895 1546 16904
rect 1492 16448 1544 16454
rect 1490 16416 1492 16425
rect 1544 16416 1546 16425
rect 1490 16351 1546 16360
rect 1688 16114 1716 16934
rect 1780 16590 1808 17478
rect 1860 16720 1912 16726
rect 1860 16662 1912 16668
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1492 15904 1544 15910
rect 1490 15872 1492 15881
rect 1676 15904 1728 15910
rect 1544 15872 1546 15881
rect 1676 15846 1728 15852
rect 1490 15807 1546 15816
rect 1492 15360 1544 15366
rect 1490 15328 1492 15337
rect 1544 15328 1546 15337
rect 1490 15263 1546 15272
rect 1492 14816 1544 14822
rect 1490 14784 1492 14793
rect 1544 14784 1546 14793
rect 1490 14719 1546 14728
rect 1492 14272 1544 14278
rect 1490 14240 1492 14249
rect 1544 14240 1546 14249
rect 1490 14175 1546 14184
rect 1400 13796 1452 13802
rect 1400 13738 1452 13744
rect 1228 11750 1348 11778
rect 1124 6180 1176 6186
rect 1124 6122 1176 6128
rect 1032 5772 1084 5778
rect 1032 5714 1084 5720
rect 1136 4554 1164 6122
rect 1228 4826 1256 11750
rect 1412 9042 1440 13738
rect 1492 13728 1544 13734
rect 1490 13696 1492 13705
rect 1544 13696 1546 13705
rect 1490 13631 1546 13640
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1504 13025 1532 13126
rect 1490 13016 1546 13025
rect 1490 12951 1546 12960
rect 1688 12850 1716 15846
rect 1872 15026 1900 16662
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12481 1532 12582
rect 1490 12472 1546 12481
rect 1490 12407 1546 12416
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11937 1532 12038
rect 1490 11928 1546 11937
rect 1490 11863 1546 11872
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1504 11393 1532 11494
rect 1490 11384 1546 11393
rect 1490 11319 1546 11328
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10849 1532 10950
rect 1490 10840 1546 10849
rect 1490 10775 1546 10784
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1504 10305 1532 10406
rect 1490 10296 1546 10305
rect 1490 10231 1546 10240
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 9761 1532 9862
rect 1490 9752 1546 9761
rect 1490 9687 1546 9696
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1412 8129 1440 8774
rect 1504 8673 1532 9318
rect 1490 8664 1546 8673
rect 1490 8599 1546 8608
rect 1596 8566 1624 12378
rect 1780 10062 1808 14758
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1688 9178 1716 9522
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1688 8498 1716 8774
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1398 8120 1454 8129
rect 1398 8055 1454 8064
rect 1308 7744 1360 7750
rect 1308 7686 1360 7692
rect 1320 6361 1348 7686
rect 1504 7585 1532 8298
rect 1490 7576 1546 7585
rect 1490 7511 1546 7520
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1306 6352 1362 6361
rect 1306 6287 1362 6296
rect 1504 5817 1532 6598
rect 1490 5808 1546 5817
rect 1490 5743 1546 5752
rect 1688 5710 1716 8298
rect 1964 7546 1992 17818
rect 2056 15570 2084 19382
rect 2332 18290 2360 27406
rect 2516 25480 2544 27474
rect 2582 26684 2890 26704
rect 2582 26682 2588 26684
rect 2644 26682 2668 26684
rect 2724 26682 2748 26684
rect 2804 26682 2828 26684
rect 2884 26682 2890 26684
rect 2644 26630 2646 26682
rect 2826 26630 2828 26682
rect 2582 26628 2588 26630
rect 2644 26628 2668 26630
rect 2724 26628 2748 26630
rect 2804 26628 2828 26630
rect 2884 26628 2890 26630
rect 2582 26608 2890 26628
rect 2582 25596 2890 25616
rect 2582 25594 2588 25596
rect 2644 25594 2668 25596
rect 2724 25594 2748 25596
rect 2804 25594 2828 25596
rect 2884 25594 2890 25596
rect 2644 25542 2646 25594
rect 2826 25542 2828 25594
rect 2582 25540 2588 25542
rect 2644 25540 2668 25542
rect 2724 25540 2748 25542
rect 2804 25540 2828 25542
rect 2884 25540 2890 25542
rect 2582 25520 2890 25540
rect 2516 25452 2636 25480
rect 2608 24818 2636 25452
rect 2596 24812 2648 24818
rect 2596 24754 2648 24760
rect 2964 24744 3016 24750
rect 2964 24686 3016 24692
rect 2504 24608 2556 24614
rect 2504 24550 2556 24556
rect 2412 20868 2464 20874
rect 2412 20810 2464 20816
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2240 17678 2268 18158
rect 2320 18148 2372 18154
rect 2320 18090 2372 18096
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2240 17202 2268 17614
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2240 16658 2268 17138
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 2148 15026 2176 15438
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2148 14414 2176 14962
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 2148 9586 2176 14214
rect 2240 11150 2268 15302
rect 2332 14414 2360 18090
rect 2424 16590 2452 20810
rect 2516 17746 2544 24550
rect 2582 24508 2890 24528
rect 2582 24506 2588 24508
rect 2644 24506 2668 24508
rect 2724 24506 2748 24508
rect 2804 24506 2828 24508
rect 2884 24506 2890 24508
rect 2644 24454 2646 24506
rect 2826 24454 2828 24506
rect 2582 24452 2588 24454
rect 2644 24452 2668 24454
rect 2724 24452 2748 24454
rect 2804 24452 2828 24454
rect 2884 24452 2890 24454
rect 2582 24432 2890 24452
rect 2976 24290 3004 24686
rect 2884 24262 3004 24290
rect 2884 24138 2912 24262
rect 2872 24132 2924 24138
rect 2872 24074 2924 24080
rect 2884 23730 2912 24074
rect 3068 23730 3096 37130
rect 3148 32428 3200 32434
rect 3148 32370 3200 32376
rect 3160 31958 3188 32370
rect 3148 31952 3200 31958
rect 3148 31894 3200 31900
rect 3252 31754 3280 45047
rect 3332 43308 3384 43314
rect 3332 43250 3384 43256
rect 3344 36582 3372 43250
rect 3332 36576 3384 36582
rect 3332 36518 3384 36524
rect 3148 31748 3200 31754
rect 3252 31726 3372 31754
rect 3148 31690 3200 31696
rect 3160 31482 3188 31690
rect 3148 31476 3200 31482
rect 3148 31418 3200 31424
rect 3148 31340 3200 31346
rect 3148 31282 3200 31288
rect 3160 30054 3188 31282
rect 3344 31226 3372 31726
rect 3252 31198 3372 31226
rect 3148 30048 3200 30054
rect 3148 29990 3200 29996
rect 3252 27606 3280 31198
rect 3332 31136 3384 31142
rect 3332 31078 3384 31084
rect 3240 27600 3292 27606
rect 3240 27542 3292 27548
rect 3344 24818 3372 31078
rect 3436 29102 3464 50186
rect 3528 49842 3556 50759
rect 3516 49836 3568 49842
rect 3516 49778 3568 49784
rect 3516 48748 3568 48754
rect 3516 48690 3568 48696
rect 3528 46102 3556 48690
rect 3712 48657 3740 52414
rect 3804 48890 3832 52550
rect 3792 48884 3844 48890
rect 3792 48826 3844 48832
rect 3698 48648 3754 48657
rect 3698 48583 3754 48592
rect 3792 48544 3844 48550
rect 3792 48486 3844 48492
rect 3698 48376 3754 48385
rect 3698 48311 3754 48320
rect 3608 47592 3660 47598
rect 3608 47534 3660 47540
rect 3620 46345 3648 47534
rect 3606 46336 3662 46345
rect 3606 46271 3662 46280
rect 3712 46186 3740 48311
rect 3620 46158 3740 46186
rect 3516 46096 3568 46102
rect 3516 46038 3568 46044
rect 3516 45960 3568 45966
rect 3516 45902 3568 45908
rect 3528 44742 3556 45902
rect 3516 44736 3568 44742
rect 3516 44678 3568 44684
rect 3516 43104 3568 43110
rect 3516 43046 3568 43052
rect 3528 41614 3556 43046
rect 3516 41608 3568 41614
rect 3516 41550 3568 41556
rect 3516 41268 3568 41274
rect 3516 41210 3568 41216
rect 3528 36666 3556 41210
rect 3620 40730 3648 46158
rect 3700 46096 3752 46102
rect 3700 46038 3752 46044
rect 3804 46050 3832 48486
rect 3896 46170 3924 56782
rect 3976 56704 4028 56710
rect 3976 56646 4028 56652
rect 3988 56409 4016 56646
rect 4080 56506 4108 66982
rect 4213 66396 4521 66416
rect 4213 66394 4219 66396
rect 4275 66394 4299 66396
rect 4355 66394 4379 66396
rect 4435 66394 4459 66396
rect 4515 66394 4521 66396
rect 4275 66342 4277 66394
rect 4457 66342 4459 66394
rect 4213 66340 4219 66342
rect 4275 66340 4299 66342
rect 4355 66340 4379 66342
rect 4435 66340 4459 66342
rect 4515 66340 4521 66342
rect 4213 66320 4521 66340
rect 4213 65308 4521 65328
rect 4213 65306 4219 65308
rect 4275 65306 4299 65308
rect 4355 65306 4379 65308
rect 4435 65306 4459 65308
rect 4515 65306 4521 65308
rect 4275 65254 4277 65306
rect 4457 65254 4459 65306
rect 4213 65252 4219 65254
rect 4275 65252 4299 65254
rect 4355 65252 4379 65254
rect 4435 65252 4459 65254
rect 4515 65252 4521 65254
rect 4213 65232 4521 65252
rect 4213 64220 4521 64240
rect 4213 64218 4219 64220
rect 4275 64218 4299 64220
rect 4355 64218 4379 64220
rect 4435 64218 4459 64220
rect 4515 64218 4521 64220
rect 4275 64166 4277 64218
rect 4457 64166 4459 64218
rect 4213 64164 4219 64166
rect 4275 64164 4299 64166
rect 4355 64164 4379 64166
rect 4435 64164 4459 64166
rect 4515 64164 4521 64166
rect 4213 64144 4521 64164
rect 4213 63132 4521 63152
rect 4213 63130 4219 63132
rect 4275 63130 4299 63132
rect 4355 63130 4379 63132
rect 4435 63130 4459 63132
rect 4515 63130 4521 63132
rect 4275 63078 4277 63130
rect 4457 63078 4459 63130
rect 4213 63076 4219 63078
rect 4275 63076 4299 63078
rect 4355 63076 4379 63078
rect 4435 63076 4459 63078
rect 4515 63076 4521 63078
rect 4213 63056 4521 63076
rect 4213 62044 4521 62064
rect 4213 62042 4219 62044
rect 4275 62042 4299 62044
rect 4355 62042 4379 62044
rect 4435 62042 4459 62044
rect 4515 62042 4521 62044
rect 4275 61990 4277 62042
rect 4457 61990 4459 62042
rect 4213 61988 4219 61990
rect 4275 61988 4299 61990
rect 4355 61988 4379 61990
rect 4435 61988 4459 61990
rect 4515 61988 4521 61990
rect 4213 61968 4521 61988
rect 4213 60956 4521 60976
rect 4213 60954 4219 60956
rect 4275 60954 4299 60956
rect 4355 60954 4379 60956
rect 4435 60954 4459 60956
rect 4515 60954 4521 60956
rect 4275 60902 4277 60954
rect 4457 60902 4459 60954
rect 4213 60900 4219 60902
rect 4275 60900 4299 60902
rect 4355 60900 4379 60902
rect 4435 60900 4459 60902
rect 4515 60900 4521 60902
rect 4213 60880 4521 60900
rect 4213 59868 4521 59888
rect 4213 59866 4219 59868
rect 4275 59866 4299 59868
rect 4355 59866 4379 59868
rect 4435 59866 4459 59868
rect 4515 59866 4521 59868
rect 4275 59814 4277 59866
rect 4457 59814 4459 59866
rect 4213 59812 4219 59814
rect 4275 59812 4299 59814
rect 4355 59812 4379 59814
rect 4435 59812 4459 59814
rect 4515 59812 4521 59814
rect 4213 59792 4521 59812
rect 4213 58780 4521 58800
rect 4213 58778 4219 58780
rect 4275 58778 4299 58780
rect 4355 58778 4379 58780
rect 4435 58778 4459 58780
rect 4515 58778 4521 58780
rect 4275 58726 4277 58778
rect 4457 58726 4459 58778
rect 4213 58724 4219 58726
rect 4275 58724 4299 58726
rect 4355 58724 4379 58726
rect 4435 58724 4459 58726
rect 4515 58724 4521 58726
rect 4213 58704 4521 58724
rect 4213 57692 4521 57712
rect 4213 57690 4219 57692
rect 4275 57690 4299 57692
rect 4355 57690 4379 57692
rect 4435 57690 4459 57692
rect 4515 57690 4521 57692
rect 4275 57638 4277 57690
rect 4457 57638 4459 57690
rect 4213 57636 4219 57638
rect 4275 57636 4299 57638
rect 4355 57636 4379 57638
rect 4435 57636 4459 57638
rect 4515 57636 4521 57638
rect 4213 57616 4521 57636
rect 4213 56604 4521 56624
rect 4213 56602 4219 56604
rect 4275 56602 4299 56604
rect 4355 56602 4379 56604
rect 4435 56602 4459 56604
rect 4515 56602 4521 56604
rect 4275 56550 4277 56602
rect 4457 56550 4459 56602
rect 4213 56548 4219 56550
rect 4275 56548 4299 56550
rect 4355 56548 4379 56550
rect 4435 56548 4459 56550
rect 4515 56548 4521 56550
rect 4213 56528 4521 56548
rect 4068 56500 4120 56506
rect 4068 56442 4120 56448
rect 3974 56400 4030 56409
rect 3974 56335 4030 56344
rect 3976 56296 4028 56302
rect 3976 56238 4028 56244
rect 3988 55706 4016 56238
rect 4080 55826 4108 56442
rect 4068 55820 4120 55826
rect 4068 55762 4120 55768
rect 3988 55678 4108 55706
rect 3976 55616 4028 55622
rect 3976 55558 4028 55564
rect 3988 55321 4016 55558
rect 3974 55312 4030 55321
rect 3974 55247 4030 55256
rect 3976 54188 4028 54194
rect 3976 54130 4028 54136
rect 3988 51097 4016 54130
rect 4080 52358 4108 55678
rect 4213 55516 4521 55536
rect 4213 55514 4219 55516
rect 4275 55514 4299 55516
rect 4355 55514 4379 55516
rect 4435 55514 4459 55516
rect 4515 55514 4521 55516
rect 4275 55462 4277 55514
rect 4457 55462 4459 55514
rect 4213 55460 4219 55462
rect 4275 55460 4299 55462
rect 4355 55460 4379 55462
rect 4435 55460 4459 55462
rect 4515 55460 4521 55462
rect 4213 55440 4521 55460
rect 4213 54428 4521 54448
rect 4213 54426 4219 54428
rect 4275 54426 4299 54428
rect 4355 54426 4379 54428
rect 4435 54426 4459 54428
rect 4515 54426 4521 54428
rect 4275 54374 4277 54426
rect 4457 54374 4459 54426
rect 4213 54372 4219 54374
rect 4275 54372 4299 54374
rect 4355 54372 4379 54374
rect 4435 54372 4459 54374
rect 4515 54372 4521 54374
rect 4213 54352 4521 54372
rect 4213 53340 4521 53360
rect 4213 53338 4219 53340
rect 4275 53338 4299 53340
rect 4355 53338 4379 53340
rect 4435 53338 4459 53340
rect 4515 53338 4521 53340
rect 4275 53286 4277 53338
rect 4457 53286 4459 53338
rect 4213 53284 4219 53286
rect 4275 53284 4299 53286
rect 4355 53284 4379 53286
rect 4435 53284 4459 53286
rect 4515 53284 4521 53286
rect 4213 53264 4521 53284
rect 4068 52352 4120 52358
rect 4068 52294 4120 52300
rect 4213 52252 4521 52272
rect 4213 52250 4219 52252
rect 4275 52250 4299 52252
rect 4355 52250 4379 52252
rect 4435 52250 4459 52252
rect 4515 52250 4521 52252
rect 4275 52198 4277 52250
rect 4457 52198 4459 52250
rect 4213 52196 4219 52198
rect 4275 52196 4299 52198
rect 4355 52196 4379 52198
rect 4435 52196 4459 52198
rect 4515 52196 4521 52198
rect 4213 52176 4521 52196
rect 4068 52012 4120 52018
rect 4068 51954 4120 51960
rect 3974 51088 4030 51097
rect 3974 51023 4030 51032
rect 3976 50924 4028 50930
rect 3976 50866 4028 50872
rect 3988 50182 4016 50866
rect 4080 50726 4108 51954
rect 4213 51164 4521 51184
rect 4213 51162 4219 51164
rect 4275 51162 4299 51164
rect 4355 51162 4379 51164
rect 4435 51162 4459 51164
rect 4515 51162 4521 51164
rect 4275 51110 4277 51162
rect 4457 51110 4459 51162
rect 4213 51108 4219 51110
rect 4275 51108 4299 51110
rect 4355 51108 4379 51110
rect 4435 51108 4459 51110
rect 4515 51108 4521 51110
rect 4213 51088 4521 51108
rect 4068 50720 4120 50726
rect 4068 50662 4120 50668
rect 4160 50720 4212 50726
rect 4160 50662 4212 50668
rect 3976 50176 4028 50182
rect 3976 50118 4028 50124
rect 3976 49836 4028 49842
rect 3976 49778 4028 49784
rect 3988 47161 4016 49778
rect 4080 49774 4108 50662
rect 4172 50386 4200 50662
rect 4160 50380 4212 50386
rect 4160 50322 4212 50328
rect 4213 50076 4521 50096
rect 4213 50074 4219 50076
rect 4275 50074 4299 50076
rect 4355 50074 4379 50076
rect 4435 50074 4459 50076
rect 4515 50074 4521 50076
rect 4275 50022 4277 50074
rect 4457 50022 4459 50074
rect 4213 50020 4219 50022
rect 4275 50020 4299 50022
rect 4355 50020 4379 50022
rect 4435 50020 4459 50022
rect 4515 50020 4521 50022
rect 4213 50000 4521 50020
rect 4068 49768 4120 49774
rect 4068 49710 4120 49716
rect 4252 49632 4304 49638
rect 4252 49574 4304 49580
rect 4264 49230 4292 49574
rect 4252 49224 4304 49230
rect 4252 49166 4304 49172
rect 4213 48988 4521 49008
rect 4213 48986 4219 48988
rect 4275 48986 4299 48988
rect 4355 48986 4379 48988
rect 4435 48986 4459 48988
rect 4515 48986 4521 48988
rect 4275 48934 4277 48986
rect 4457 48934 4459 48986
rect 4213 48932 4219 48934
rect 4275 48932 4299 48934
rect 4355 48932 4379 48934
rect 4435 48932 4459 48934
rect 4515 48932 4521 48934
rect 4213 48912 4521 48932
rect 4213 47900 4521 47920
rect 4213 47898 4219 47900
rect 4275 47898 4299 47900
rect 4355 47898 4379 47900
rect 4435 47898 4459 47900
rect 4515 47898 4521 47900
rect 4275 47846 4277 47898
rect 4457 47846 4459 47898
rect 4213 47844 4219 47846
rect 4275 47844 4299 47846
rect 4355 47844 4379 47846
rect 4435 47844 4459 47846
rect 4515 47844 4521 47846
rect 4213 47824 4521 47844
rect 4160 47456 4212 47462
rect 4160 47398 4212 47404
rect 3974 47152 4030 47161
rect 3974 47087 4030 47096
rect 4172 47002 4200 47398
rect 3988 46974 4200 47002
rect 3988 46646 4016 46974
rect 4068 46912 4120 46918
rect 4068 46854 4120 46860
rect 3976 46640 4028 46646
rect 3976 46582 4028 46588
rect 3976 46436 4028 46442
rect 3976 46378 4028 46384
rect 3884 46164 3936 46170
rect 3884 46106 3936 46112
rect 3608 40724 3660 40730
rect 3608 40666 3660 40672
rect 3608 38208 3660 38214
rect 3608 38150 3660 38156
rect 3620 36802 3648 38150
rect 3712 36922 3740 46038
rect 3804 46022 3924 46050
rect 3988 46034 4016 46378
rect 3792 45892 3844 45898
rect 3792 45834 3844 45840
rect 3804 44878 3832 45834
rect 3792 44872 3844 44878
rect 3792 44814 3844 44820
rect 3792 44736 3844 44742
rect 3792 44678 3844 44684
rect 3804 38554 3832 44678
rect 3896 41206 3924 46022
rect 3976 46028 4028 46034
rect 3976 45970 4028 45976
rect 4080 45966 4108 46854
rect 4213 46812 4521 46832
rect 4213 46810 4219 46812
rect 4275 46810 4299 46812
rect 4355 46810 4379 46812
rect 4435 46810 4459 46812
rect 4515 46810 4521 46812
rect 4275 46758 4277 46810
rect 4457 46758 4459 46810
rect 4213 46756 4219 46758
rect 4275 46756 4299 46758
rect 4355 46756 4379 46758
rect 4435 46756 4459 46758
rect 4515 46756 4521 46758
rect 4213 46736 4521 46756
rect 4068 45960 4120 45966
rect 4068 45902 4120 45908
rect 3976 45824 4028 45830
rect 3976 45766 4028 45772
rect 3988 45286 4016 45766
rect 4213 45724 4521 45744
rect 4213 45722 4219 45724
rect 4275 45722 4299 45724
rect 4355 45722 4379 45724
rect 4435 45722 4459 45724
rect 4515 45722 4521 45724
rect 4275 45670 4277 45722
rect 4457 45670 4459 45722
rect 4213 45668 4219 45670
rect 4275 45668 4299 45670
rect 4355 45668 4379 45670
rect 4435 45668 4459 45670
rect 4515 45668 4521 45670
rect 4213 45648 4521 45668
rect 4068 45416 4120 45422
rect 4068 45358 4120 45364
rect 3976 45280 4028 45286
rect 3976 45222 4028 45228
rect 3974 45112 4030 45121
rect 3974 45047 4030 45056
rect 3988 42702 4016 45047
rect 4080 42770 4108 45358
rect 4213 44636 4521 44656
rect 4213 44634 4219 44636
rect 4275 44634 4299 44636
rect 4355 44634 4379 44636
rect 4435 44634 4459 44636
rect 4515 44634 4521 44636
rect 4275 44582 4277 44634
rect 4457 44582 4459 44634
rect 4213 44580 4219 44582
rect 4275 44580 4299 44582
rect 4355 44580 4379 44582
rect 4435 44580 4459 44582
rect 4515 44580 4521 44582
rect 4213 44560 4521 44580
rect 4213 43548 4521 43568
rect 4213 43546 4219 43548
rect 4275 43546 4299 43548
rect 4355 43546 4379 43548
rect 4435 43546 4459 43548
rect 4515 43546 4521 43548
rect 4275 43494 4277 43546
rect 4457 43494 4459 43546
rect 4213 43492 4219 43494
rect 4275 43492 4299 43494
rect 4355 43492 4379 43494
rect 4435 43492 4459 43494
rect 4515 43492 4521 43494
rect 4213 43472 4521 43492
rect 4068 42764 4120 42770
rect 4068 42706 4120 42712
rect 3976 42696 4028 42702
rect 3976 42638 4028 42644
rect 3976 42016 4028 42022
rect 3976 41958 4028 41964
rect 3884 41200 3936 41206
rect 3884 41142 3936 41148
rect 3988 41138 4016 41958
rect 4080 41857 4108 42706
rect 4213 42460 4521 42480
rect 4213 42458 4219 42460
rect 4275 42458 4299 42460
rect 4355 42458 4379 42460
rect 4435 42458 4459 42460
rect 4515 42458 4521 42460
rect 4275 42406 4277 42458
rect 4457 42406 4459 42458
rect 4213 42404 4219 42406
rect 4275 42404 4299 42406
rect 4355 42404 4379 42406
rect 4435 42404 4459 42406
rect 4515 42404 4521 42406
rect 4213 42384 4521 42404
rect 4066 41848 4122 41857
rect 4066 41783 4122 41792
rect 4068 41744 4120 41750
rect 4068 41686 4120 41692
rect 4080 41256 4108 41686
rect 4158 41576 4214 41585
rect 4158 41511 4160 41520
rect 4212 41511 4214 41520
rect 4160 41482 4212 41488
rect 4213 41372 4521 41392
rect 4213 41370 4219 41372
rect 4275 41370 4299 41372
rect 4355 41370 4379 41372
rect 4435 41370 4459 41372
rect 4515 41370 4521 41372
rect 4275 41318 4277 41370
rect 4457 41318 4459 41370
rect 4213 41316 4219 41318
rect 4275 41316 4299 41318
rect 4355 41316 4379 41318
rect 4435 41316 4459 41318
rect 4515 41316 4521 41318
rect 4213 41296 4521 41316
rect 4080 41228 4200 41256
rect 3976 41132 4028 41138
rect 3976 41074 4028 41080
rect 3884 40996 3936 41002
rect 3884 40938 3936 40944
rect 3896 39794 3924 40938
rect 3988 40186 4016 41074
rect 4172 40372 4200 41228
rect 4526 41168 4582 41177
rect 4526 41103 4582 41112
rect 4436 40928 4488 40934
rect 4436 40870 4488 40876
rect 4448 40730 4476 40870
rect 4436 40724 4488 40730
rect 4436 40666 4488 40672
rect 4540 40508 4568 41103
rect 4632 40662 4660 71674
rect 4724 55214 4752 73782
rect 4816 73778 4844 74190
rect 4988 74180 5040 74186
rect 4988 74122 5040 74128
rect 5000 73778 5028 74122
rect 4804 73772 4856 73778
rect 4804 73714 4856 73720
rect 4988 73772 5040 73778
rect 4988 73714 5040 73720
rect 4988 73636 5040 73642
rect 4988 73578 5040 73584
rect 4804 73364 4856 73370
rect 4804 73306 4856 73312
rect 4712 55208 4764 55214
rect 4712 55150 4764 55156
rect 4712 49972 4764 49978
rect 4712 49914 4764 49920
rect 4620 40656 4672 40662
rect 4620 40598 4672 40604
rect 4540 40480 4660 40508
rect 4080 40344 4200 40372
rect 3976 40180 4028 40186
rect 3976 40122 4028 40128
rect 3896 39766 4016 39794
rect 3884 38888 3936 38894
rect 3884 38830 3936 38836
rect 3792 38548 3844 38554
rect 3792 38490 3844 38496
rect 3896 37670 3924 38830
rect 3884 37664 3936 37670
rect 3884 37606 3936 37612
rect 3700 36916 3752 36922
rect 3700 36858 3752 36864
rect 3792 36848 3844 36854
rect 3620 36774 3740 36802
rect 3792 36790 3844 36796
rect 3528 36638 3648 36666
rect 3516 36576 3568 36582
rect 3516 36518 3568 36524
rect 3424 29096 3476 29102
rect 3424 29038 3476 29044
rect 3424 28960 3476 28966
rect 3424 28902 3476 28908
rect 3436 28098 3464 28902
rect 3528 28218 3556 36518
rect 3620 36378 3648 36638
rect 3608 36372 3660 36378
rect 3608 36314 3660 36320
rect 3712 31754 3740 36774
rect 3804 36174 3832 36790
rect 3884 36576 3936 36582
rect 3884 36518 3936 36524
rect 3792 36168 3844 36174
rect 3792 36110 3844 36116
rect 3804 34542 3832 36110
rect 3792 34536 3844 34542
rect 3792 34478 3844 34484
rect 3620 31726 3740 31754
rect 3516 28212 3568 28218
rect 3516 28154 3568 28160
rect 3436 28070 3556 28098
rect 3424 27600 3476 27606
rect 3424 27542 3476 27548
rect 3332 24812 3384 24818
rect 3332 24754 3384 24760
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 3056 23724 3108 23730
rect 3056 23666 3108 23672
rect 2884 23610 2912 23666
rect 2884 23582 3004 23610
rect 2582 23420 2890 23440
rect 2582 23418 2588 23420
rect 2644 23418 2668 23420
rect 2724 23418 2748 23420
rect 2804 23418 2828 23420
rect 2884 23418 2890 23420
rect 2644 23366 2646 23418
rect 2826 23366 2828 23418
rect 2582 23364 2588 23366
rect 2644 23364 2668 23366
rect 2724 23364 2748 23366
rect 2804 23364 2828 23366
rect 2884 23364 2890 23366
rect 2582 23344 2890 23364
rect 2976 23050 3004 23582
rect 3332 23588 3384 23594
rect 3332 23530 3384 23536
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 2964 23044 3016 23050
rect 2964 22986 3016 22992
rect 2976 22574 3004 22986
rect 3056 22976 3108 22982
rect 3056 22918 3108 22924
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 2582 22332 2890 22352
rect 2582 22330 2588 22332
rect 2644 22330 2668 22332
rect 2724 22330 2748 22332
rect 2804 22330 2828 22332
rect 2884 22330 2890 22332
rect 2644 22278 2646 22330
rect 2826 22278 2828 22330
rect 2582 22276 2588 22278
rect 2644 22276 2668 22278
rect 2724 22276 2748 22278
rect 2804 22276 2828 22278
rect 2884 22276 2890 22278
rect 2582 22256 2890 22276
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2700 21622 2728 21966
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 2688 21616 2740 21622
rect 2688 21558 2740 21564
rect 2976 21350 3004 21898
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2582 21244 2890 21264
rect 2582 21242 2588 21244
rect 2644 21242 2668 21244
rect 2724 21242 2748 21244
rect 2804 21242 2828 21244
rect 2884 21242 2890 21244
rect 2644 21190 2646 21242
rect 2826 21190 2828 21242
rect 2582 21188 2588 21190
rect 2644 21188 2668 21190
rect 2724 21188 2748 21190
rect 2804 21188 2828 21190
rect 2884 21188 2890 21190
rect 2582 21168 2890 21188
rect 3068 20942 3096 22918
rect 3160 21554 3188 23462
rect 3240 22636 3292 22642
rect 3240 22578 3292 22584
rect 3148 21548 3200 21554
rect 3148 21490 3200 21496
rect 3252 21350 3280 22578
rect 3148 21344 3200 21350
rect 3148 21286 3200 21292
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 2582 20156 2890 20176
rect 2582 20154 2588 20156
rect 2644 20154 2668 20156
rect 2724 20154 2748 20156
rect 2804 20154 2828 20156
rect 2884 20154 2890 20156
rect 2644 20102 2646 20154
rect 2826 20102 2828 20154
rect 2582 20100 2588 20102
rect 2644 20100 2668 20102
rect 2724 20100 2748 20102
rect 2804 20100 2828 20102
rect 2884 20100 2890 20102
rect 2582 20080 2890 20100
rect 2582 19068 2890 19088
rect 2582 19066 2588 19068
rect 2644 19066 2668 19068
rect 2724 19066 2748 19068
rect 2804 19066 2828 19068
rect 2884 19066 2890 19068
rect 2644 19014 2646 19066
rect 2826 19014 2828 19066
rect 2582 19012 2588 19014
rect 2644 19012 2668 19014
rect 2724 19012 2748 19014
rect 2804 19012 2828 19014
rect 2884 19012 2890 19014
rect 2582 18992 2890 19012
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2582 17980 2890 18000
rect 2582 17978 2588 17980
rect 2644 17978 2668 17980
rect 2724 17978 2748 17980
rect 2804 17978 2828 17980
rect 2884 17978 2890 17980
rect 2644 17926 2646 17978
rect 2826 17926 2828 17978
rect 2582 17924 2588 17926
rect 2644 17924 2668 17926
rect 2724 17924 2748 17926
rect 2804 17924 2828 17926
rect 2884 17924 2890 17926
rect 2582 17904 2890 17924
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 2582 16892 2890 16912
rect 2582 16890 2588 16892
rect 2644 16890 2668 16892
rect 2724 16890 2748 16892
rect 2804 16890 2828 16892
rect 2884 16890 2890 16892
rect 2644 16838 2646 16890
rect 2826 16838 2828 16890
rect 2582 16836 2588 16838
rect 2644 16836 2668 16838
rect 2724 16836 2748 16838
rect 2804 16836 2828 16838
rect 2884 16836 2890 16838
rect 2582 16816 2890 16836
rect 2976 16726 3004 18022
rect 2964 16720 3016 16726
rect 2964 16662 3016 16668
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2582 15804 2890 15824
rect 2582 15802 2588 15804
rect 2644 15802 2668 15804
rect 2724 15802 2748 15804
rect 2804 15802 2828 15804
rect 2884 15802 2890 15804
rect 2644 15750 2646 15802
rect 2826 15750 2828 15802
rect 2582 15748 2588 15750
rect 2644 15748 2668 15750
rect 2724 15748 2748 15750
rect 2804 15748 2828 15750
rect 2884 15748 2890 15750
rect 2582 15728 2890 15748
rect 2976 15638 3004 16390
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2964 15632 3016 15638
rect 2964 15574 3016 15580
rect 3068 14906 3096 15846
rect 2976 14878 3096 14906
rect 2582 14716 2890 14736
rect 2582 14714 2588 14716
rect 2644 14714 2668 14716
rect 2724 14714 2748 14716
rect 2804 14714 2828 14716
rect 2884 14714 2890 14716
rect 2644 14662 2646 14714
rect 2826 14662 2828 14714
rect 2582 14660 2588 14662
rect 2644 14660 2668 14662
rect 2724 14660 2748 14662
rect 2804 14660 2828 14662
rect 2884 14660 2890 14662
rect 2582 14640 2890 14660
rect 2976 14550 3004 14878
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 2964 14544 3016 14550
rect 2964 14486 3016 14492
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2516 13530 2544 14350
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2582 13628 2890 13648
rect 2582 13626 2588 13628
rect 2644 13626 2668 13628
rect 2724 13626 2748 13628
rect 2804 13626 2828 13628
rect 2884 13626 2890 13628
rect 2644 13574 2646 13626
rect 2826 13574 2828 13626
rect 2582 13572 2588 13574
rect 2644 13572 2668 13574
rect 2724 13572 2748 13574
rect 2804 13572 2828 13574
rect 2884 13572 2890 13574
rect 2582 13552 2890 13572
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2792 12850 2820 13262
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2582 12540 2890 12560
rect 2582 12538 2588 12540
rect 2644 12538 2668 12540
rect 2724 12538 2748 12540
rect 2804 12538 2828 12540
rect 2884 12538 2890 12540
rect 2644 12486 2646 12538
rect 2826 12486 2828 12538
rect 2582 12484 2588 12486
rect 2644 12484 2668 12486
rect 2724 12484 2748 12486
rect 2804 12484 2828 12486
rect 2884 12484 2890 12486
rect 2582 12464 2890 12484
rect 2582 11452 2890 11472
rect 2582 11450 2588 11452
rect 2644 11450 2668 11452
rect 2724 11450 2748 11452
rect 2804 11450 2828 11452
rect 2884 11450 2890 11452
rect 2644 11398 2646 11450
rect 2826 11398 2828 11450
rect 2582 11396 2588 11398
rect 2644 11396 2668 11398
rect 2724 11396 2748 11398
rect 2804 11396 2828 11398
rect 2884 11396 2890 11398
rect 2582 11376 2890 11396
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2976 10674 3004 14214
rect 3068 11762 3096 14758
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2582 10364 2890 10384
rect 2582 10362 2588 10364
rect 2644 10362 2668 10364
rect 2724 10362 2748 10364
rect 2804 10362 2828 10364
rect 2884 10362 2890 10364
rect 2644 10310 2646 10362
rect 2826 10310 2828 10362
rect 2582 10308 2588 10310
rect 2644 10308 2668 10310
rect 2724 10308 2748 10310
rect 2804 10308 2828 10310
rect 2884 10308 2890 10310
rect 2582 10288 2890 10308
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2332 9217 2360 9318
rect 2582 9276 2890 9296
rect 2582 9274 2588 9276
rect 2644 9274 2668 9276
rect 2724 9274 2748 9276
rect 2804 9274 2828 9276
rect 2884 9274 2890 9276
rect 2644 9222 2646 9274
rect 2826 9222 2828 9274
rect 2582 9220 2588 9222
rect 2644 9220 2668 9222
rect 2724 9220 2748 9222
rect 2804 9220 2828 9222
rect 2884 9220 2890 9222
rect 2318 9208 2374 9217
rect 2582 9200 2890 9220
rect 2318 9143 2374 9152
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2240 8634 2268 8910
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2148 7886 2176 8434
rect 2332 7886 2360 9046
rect 3068 8974 3096 9998
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3068 8566 3096 8910
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2582 8188 2890 8208
rect 2582 8186 2588 8188
rect 2644 8186 2668 8188
rect 2724 8186 2748 8188
rect 2804 8186 2828 8188
rect 2884 8186 2890 8188
rect 2644 8134 2646 8186
rect 2826 8134 2828 8186
rect 2582 8132 2588 8134
rect 2644 8132 2668 8134
rect 2724 8132 2748 8134
rect 2804 8132 2828 8134
rect 2884 8132 2890 8134
rect 2582 8112 2890 8132
rect 2976 8022 3004 8230
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1504 5273 1532 5510
rect 1490 5264 1546 5273
rect 1490 5199 1546 5208
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1216 4820 1268 4826
rect 1216 4762 1268 4768
rect 1504 4729 1532 4966
rect 1490 4720 1546 4729
rect 1490 4655 1546 4664
rect 1124 4548 1176 4554
rect 1124 4490 1176 4496
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1504 4185 1532 4422
rect 1490 4176 1546 4185
rect 1490 4111 1546 4120
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1412 2553 1440 3334
rect 1504 3097 1532 3878
rect 1688 3534 1716 4422
rect 1964 3534 1992 7346
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2056 7041 2084 7142
rect 2042 7032 2098 7041
rect 2042 6967 2098 6976
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2056 5302 2084 5646
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1490 3088 1546 3097
rect 1490 3023 1546 3032
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1398 2544 1454 2553
rect 1398 2479 1454 2488
rect 1400 2304 1452 2310
rect 1400 2246 1452 2252
rect 1412 921 1440 2246
rect 1504 2009 1532 2790
rect 1688 2446 1716 3334
rect 2148 2446 2176 5510
rect 2240 4146 2268 7686
rect 2332 6458 2360 7822
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 2582 7100 2890 7120
rect 2582 7098 2588 7100
rect 2644 7098 2668 7100
rect 2724 7098 2748 7100
rect 2804 7098 2828 7100
rect 2884 7098 2890 7100
rect 2644 7046 2646 7098
rect 2826 7046 2828 7098
rect 2582 7044 2588 7046
rect 2644 7044 2668 7046
rect 2724 7044 2748 7046
rect 2804 7044 2828 7046
rect 2884 7044 2890 7046
rect 2582 7024 2890 7044
rect 2976 6866 3004 7686
rect 3068 7410 3096 7686
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3160 6866 3188 21286
rect 3344 19378 3372 23530
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3252 15570 3280 15982
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 12238 3280 15302
rect 3344 15026 3372 17274
rect 3436 16574 3464 27542
rect 3528 21434 3556 28070
rect 3620 23730 3648 31726
rect 3896 28762 3924 36518
rect 3988 36394 4016 39766
rect 4080 36582 4108 40344
rect 4213 40284 4521 40304
rect 4213 40282 4219 40284
rect 4275 40282 4299 40284
rect 4355 40282 4379 40284
rect 4435 40282 4459 40284
rect 4515 40282 4521 40284
rect 4275 40230 4277 40282
rect 4457 40230 4459 40282
rect 4213 40228 4219 40230
rect 4275 40228 4299 40230
rect 4355 40228 4379 40230
rect 4435 40228 4459 40230
rect 4515 40228 4521 40230
rect 4213 40208 4521 40228
rect 4213 39196 4521 39216
rect 4213 39194 4219 39196
rect 4275 39194 4299 39196
rect 4355 39194 4379 39196
rect 4435 39194 4459 39196
rect 4515 39194 4521 39196
rect 4275 39142 4277 39194
rect 4457 39142 4459 39194
rect 4213 39140 4219 39142
rect 4275 39140 4299 39142
rect 4355 39140 4379 39142
rect 4435 39140 4459 39142
rect 4515 39140 4521 39142
rect 4213 39120 4521 39140
rect 4213 38108 4521 38128
rect 4213 38106 4219 38108
rect 4275 38106 4299 38108
rect 4355 38106 4379 38108
rect 4435 38106 4459 38108
rect 4515 38106 4521 38108
rect 4275 38054 4277 38106
rect 4457 38054 4459 38106
rect 4213 38052 4219 38054
rect 4275 38052 4299 38054
rect 4355 38052 4379 38054
rect 4435 38052 4459 38054
rect 4515 38052 4521 38054
rect 4213 38032 4521 38052
rect 4213 37020 4521 37040
rect 4213 37018 4219 37020
rect 4275 37018 4299 37020
rect 4355 37018 4379 37020
rect 4435 37018 4459 37020
rect 4515 37018 4521 37020
rect 4275 36966 4277 37018
rect 4457 36966 4459 37018
rect 4213 36964 4219 36966
rect 4275 36964 4299 36966
rect 4355 36964 4379 36966
rect 4435 36964 4459 36966
rect 4515 36964 4521 36966
rect 4213 36944 4521 36964
rect 4068 36576 4120 36582
rect 4068 36518 4120 36524
rect 4344 36576 4396 36582
rect 4344 36518 4396 36524
rect 3988 36366 4108 36394
rect 3976 35216 4028 35222
rect 3976 35158 4028 35164
rect 3884 28756 3936 28762
rect 3884 28698 3936 28704
rect 3884 28212 3936 28218
rect 3884 28154 3936 28160
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3608 23724 3660 23730
rect 3608 23666 3660 23672
rect 3608 22024 3660 22030
rect 3608 21966 3660 21972
rect 3620 21690 3648 21966
rect 3608 21684 3660 21690
rect 3608 21626 3660 21632
rect 3712 21570 3740 24550
rect 3792 23656 3844 23662
rect 3792 23598 3844 23604
rect 3804 23118 3832 23598
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 3804 21962 3832 23054
rect 3792 21956 3844 21962
rect 3792 21898 3844 21904
rect 3712 21542 3832 21570
rect 3528 21406 3740 21434
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3436 16546 3556 16574
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3436 15026 3464 15506
rect 3528 15094 3556 16546
rect 3516 15088 3568 15094
rect 3516 15030 3568 15036
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 3436 14906 3464 14962
rect 3344 14878 3464 14906
rect 3344 14414 3372 14878
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3344 13870 3372 14350
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3436 13462 3464 14758
rect 3620 13870 3648 21286
rect 3712 16114 3740 21406
rect 3804 18358 3832 21542
rect 3792 18352 3844 18358
rect 3792 18294 3844 18300
rect 3792 16788 3844 16794
rect 3792 16730 3844 16736
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3620 13326 3648 13806
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3344 8974 3372 12718
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3252 7410 3280 7754
rect 3436 7410 3464 11018
rect 3620 10130 3648 13262
rect 3804 12850 3832 16730
rect 3896 14414 3924 28154
rect 3988 23118 4016 35158
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3988 21622 4016 21830
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 4080 17882 4108 36366
rect 4356 36174 4384 36518
rect 4344 36168 4396 36174
rect 4344 36110 4396 36116
rect 4213 35932 4521 35952
rect 4213 35930 4219 35932
rect 4275 35930 4299 35932
rect 4355 35930 4379 35932
rect 4435 35930 4459 35932
rect 4515 35930 4521 35932
rect 4275 35878 4277 35930
rect 4457 35878 4459 35930
rect 4213 35876 4219 35878
rect 4275 35876 4299 35878
rect 4355 35876 4379 35878
rect 4435 35876 4459 35878
rect 4515 35876 4521 35878
rect 4213 35856 4521 35876
rect 4252 35760 4304 35766
rect 4252 35702 4304 35708
rect 4264 35018 4292 35702
rect 4632 35630 4660 40480
rect 4620 35624 4672 35630
rect 4620 35566 4672 35572
rect 4252 35012 4304 35018
rect 4252 34954 4304 34960
rect 4213 34844 4521 34864
rect 4213 34842 4219 34844
rect 4275 34842 4299 34844
rect 4355 34842 4379 34844
rect 4435 34842 4459 34844
rect 4515 34842 4521 34844
rect 4275 34790 4277 34842
rect 4457 34790 4459 34842
rect 4213 34788 4219 34790
rect 4275 34788 4299 34790
rect 4355 34788 4379 34790
rect 4435 34788 4459 34790
rect 4515 34788 4521 34790
rect 4213 34768 4521 34788
rect 4618 34368 4674 34377
rect 4618 34303 4674 34312
rect 4213 33756 4521 33776
rect 4213 33754 4219 33756
rect 4275 33754 4299 33756
rect 4355 33754 4379 33756
rect 4435 33754 4459 33756
rect 4515 33754 4521 33756
rect 4275 33702 4277 33754
rect 4457 33702 4459 33754
rect 4213 33700 4219 33702
rect 4275 33700 4299 33702
rect 4355 33700 4379 33702
rect 4435 33700 4459 33702
rect 4515 33700 4521 33702
rect 4213 33680 4521 33700
rect 4213 32668 4521 32688
rect 4213 32666 4219 32668
rect 4275 32666 4299 32668
rect 4355 32666 4379 32668
rect 4435 32666 4459 32668
rect 4515 32666 4521 32668
rect 4275 32614 4277 32666
rect 4457 32614 4459 32666
rect 4213 32612 4219 32614
rect 4275 32612 4299 32614
rect 4355 32612 4379 32614
rect 4435 32612 4459 32614
rect 4515 32612 4521 32614
rect 4213 32592 4521 32612
rect 4213 31580 4521 31600
rect 4213 31578 4219 31580
rect 4275 31578 4299 31580
rect 4355 31578 4379 31580
rect 4435 31578 4459 31580
rect 4515 31578 4521 31580
rect 4275 31526 4277 31578
rect 4457 31526 4459 31578
rect 4213 31524 4219 31526
rect 4275 31524 4299 31526
rect 4355 31524 4379 31526
rect 4435 31524 4459 31526
rect 4515 31524 4521 31526
rect 4213 31504 4521 31524
rect 4213 30492 4521 30512
rect 4213 30490 4219 30492
rect 4275 30490 4299 30492
rect 4355 30490 4379 30492
rect 4435 30490 4459 30492
rect 4515 30490 4521 30492
rect 4275 30438 4277 30490
rect 4457 30438 4459 30490
rect 4213 30436 4219 30438
rect 4275 30436 4299 30438
rect 4355 30436 4379 30438
rect 4435 30436 4459 30438
rect 4515 30436 4521 30438
rect 4213 30416 4521 30436
rect 4213 29404 4521 29424
rect 4213 29402 4219 29404
rect 4275 29402 4299 29404
rect 4355 29402 4379 29404
rect 4435 29402 4459 29404
rect 4515 29402 4521 29404
rect 4275 29350 4277 29402
rect 4457 29350 4459 29402
rect 4213 29348 4219 29350
rect 4275 29348 4299 29350
rect 4355 29348 4379 29350
rect 4435 29348 4459 29350
rect 4515 29348 4521 29350
rect 4213 29328 4521 29348
rect 4213 28316 4521 28336
rect 4213 28314 4219 28316
rect 4275 28314 4299 28316
rect 4355 28314 4379 28316
rect 4435 28314 4459 28316
rect 4515 28314 4521 28316
rect 4275 28262 4277 28314
rect 4457 28262 4459 28314
rect 4213 28260 4219 28262
rect 4275 28260 4299 28262
rect 4355 28260 4379 28262
rect 4435 28260 4459 28262
rect 4515 28260 4521 28262
rect 4213 28240 4521 28260
rect 4632 28098 4660 34303
rect 4724 31142 4752 49914
rect 4816 36650 4844 73306
rect 5000 70394 5028 73578
rect 5000 70366 5120 70394
rect 4896 51264 4948 51270
rect 4896 51206 4948 51212
rect 4908 50930 4936 51206
rect 5092 51074 5120 70366
rect 5356 65136 5408 65142
rect 5356 65078 5408 65084
rect 5092 51046 5304 51074
rect 4896 50924 4948 50930
rect 4896 50866 4948 50872
rect 4804 36644 4856 36650
rect 4804 36586 4856 36592
rect 4804 36100 4856 36106
rect 4804 36042 4856 36048
rect 4816 34950 4844 36042
rect 4804 34944 4856 34950
rect 4804 34886 4856 34892
rect 4712 31136 4764 31142
rect 4712 31078 4764 31084
rect 4712 30932 4764 30938
rect 4712 30874 4764 30880
rect 4724 28966 4752 30874
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 4540 28070 4660 28098
rect 4540 27606 4568 28070
rect 4620 28008 4672 28014
rect 4620 27950 4672 27956
rect 4528 27600 4580 27606
rect 4528 27542 4580 27548
rect 4213 27228 4521 27248
rect 4213 27226 4219 27228
rect 4275 27226 4299 27228
rect 4355 27226 4379 27228
rect 4435 27226 4459 27228
rect 4515 27226 4521 27228
rect 4275 27174 4277 27226
rect 4457 27174 4459 27226
rect 4213 27172 4219 27174
rect 4275 27172 4299 27174
rect 4355 27172 4379 27174
rect 4435 27172 4459 27174
rect 4515 27172 4521 27174
rect 4213 27152 4521 27172
rect 4213 26140 4521 26160
rect 4213 26138 4219 26140
rect 4275 26138 4299 26140
rect 4355 26138 4379 26140
rect 4435 26138 4459 26140
rect 4515 26138 4521 26140
rect 4275 26086 4277 26138
rect 4457 26086 4459 26138
rect 4213 26084 4219 26086
rect 4275 26084 4299 26086
rect 4355 26084 4379 26086
rect 4435 26084 4459 26086
rect 4515 26084 4521 26086
rect 4213 26064 4521 26084
rect 4213 25052 4521 25072
rect 4213 25050 4219 25052
rect 4275 25050 4299 25052
rect 4355 25050 4379 25052
rect 4435 25050 4459 25052
rect 4515 25050 4521 25052
rect 4275 24998 4277 25050
rect 4457 24998 4459 25050
rect 4213 24996 4219 24998
rect 4275 24996 4299 24998
rect 4355 24996 4379 24998
rect 4435 24996 4459 24998
rect 4515 24996 4521 24998
rect 4213 24976 4521 24996
rect 4213 23964 4521 23984
rect 4213 23962 4219 23964
rect 4275 23962 4299 23964
rect 4355 23962 4379 23964
rect 4435 23962 4459 23964
rect 4515 23962 4521 23964
rect 4275 23910 4277 23962
rect 4457 23910 4459 23962
rect 4213 23908 4219 23910
rect 4275 23908 4299 23910
rect 4355 23908 4379 23910
rect 4435 23908 4459 23910
rect 4515 23908 4521 23910
rect 4213 23888 4521 23908
rect 4213 22876 4521 22896
rect 4213 22874 4219 22876
rect 4275 22874 4299 22876
rect 4355 22874 4379 22876
rect 4435 22874 4459 22876
rect 4515 22874 4521 22876
rect 4275 22822 4277 22874
rect 4457 22822 4459 22874
rect 4213 22820 4219 22822
rect 4275 22820 4299 22822
rect 4355 22820 4379 22822
rect 4435 22820 4459 22822
rect 4515 22820 4521 22822
rect 4213 22800 4521 22820
rect 4213 21788 4521 21808
rect 4213 21786 4219 21788
rect 4275 21786 4299 21788
rect 4355 21786 4379 21788
rect 4435 21786 4459 21788
rect 4515 21786 4521 21788
rect 4275 21734 4277 21786
rect 4457 21734 4459 21786
rect 4213 21732 4219 21734
rect 4275 21732 4299 21734
rect 4355 21732 4379 21734
rect 4435 21732 4459 21734
rect 4515 21732 4521 21734
rect 4213 21712 4521 21732
rect 4213 20700 4521 20720
rect 4213 20698 4219 20700
rect 4275 20698 4299 20700
rect 4355 20698 4379 20700
rect 4435 20698 4459 20700
rect 4515 20698 4521 20700
rect 4275 20646 4277 20698
rect 4457 20646 4459 20698
rect 4213 20644 4219 20646
rect 4275 20644 4299 20646
rect 4355 20644 4379 20646
rect 4435 20644 4459 20646
rect 4515 20644 4521 20646
rect 4213 20624 4521 20644
rect 4213 19612 4521 19632
rect 4213 19610 4219 19612
rect 4275 19610 4299 19612
rect 4355 19610 4379 19612
rect 4435 19610 4459 19612
rect 4515 19610 4521 19612
rect 4275 19558 4277 19610
rect 4457 19558 4459 19610
rect 4213 19556 4219 19558
rect 4275 19556 4299 19558
rect 4355 19556 4379 19558
rect 4435 19556 4459 19558
rect 4515 19556 4521 19558
rect 4213 19536 4521 19556
rect 4213 18524 4521 18544
rect 4213 18522 4219 18524
rect 4275 18522 4299 18524
rect 4355 18522 4379 18524
rect 4435 18522 4459 18524
rect 4515 18522 4521 18524
rect 4275 18470 4277 18522
rect 4457 18470 4459 18522
rect 4213 18468 4219 18470
rect 4275 18468 4299 18470
rect 4355 18468 4379 18470
rect 4435 18468 4459 18470
rect 4515 18468 4521 18470
rect 4213 18448 4521 18468
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4213 17436 4521 17456
rect 4213 17434 4219 17436
rect 4275 17434 4299 17436
rect 4355 17434 4379 17436
rect 4435 17434 4459 17436
rect 4515 17434 4521 17436
rect 4275 17382 4277 17434
rect 4457 17382 4459 17434
rect 4213 17380 4219 17382
rect 4275 17380 4299 17382
rect 4355 17380 4379 17382
rect 4435 17380 4459 17382
rect 4515 17380 4521 17382
rect 4213 17360 4521 17380
rect 4213 16348 4521 16368
rect 4213 16346 4219 16348
rect 4275 16346 4299 16348
rect 4355 16346 4379 16348
rect 4435 16346 4459 16348
rect 4515 16346 4521 16348
rect 4275 16294 4277 16346
rect 4457 16294 4459 16346
rect 4213 16292 4219 16294
rect 4275 16292 4299 16294
rect 4355 16292 4379 16294
rect 4435 16292 4459 16294
rect 4515 16292 4521 16294
rect 4213 16272 4521 16292
rect 4213 15260 4521 15280
rect 4213 15258 4219 15260
rect 4275 15258 4299 15260
rect 4355 15258 4379 15260
rect 4435 15258 4459 15260
rect 4515 15258 4521 15260
rect 4275 15206 4277 15258
rect 4457 15206 4459 15258
rect 4213 15204 4219 15206
rect 4275 15204 4299 15206
rect 4355 15204 4379 15206
rect 4435 15204 4459 15206
rect 4515 15204 4521 15206
rect 4213 15184 4521 15204
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3896 13938 3924 14214
rect 4213 14172 4521 14192
rect 4213 14170 4219 14172
rect 4275 14170 4299 14172
rect 4355 14170 4379 14172
rect 4435 14170 4459 14172
rect 4515 14170 4521 14172
rect 4275 14118 4277 14170
rect 4457 14118 4459 14170
rect 4213 14116 4219 14118
rect 4275 14116 4299 14118
rect 4355 14116 4379 14118
rect 4435 14116 4459 14118
rect 4515 14116 4521 14118
rect 4213 14096 4521 14116
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 4213 13084 4521 13104
rect 4213 13082 4219 13084
rect 4275 13082 4299 13084
rect 4355 13082 4379 13084
rect 4435 13082 4459 13084
rect 4515 13082 4521 13084
rect 4275 13030 4277 13082
rect 4457 13030 4459 13082
rect 4213 13028 4219 13030
rect 4275 13028 4299 13030
rect 4355 13028 4379 13030
rect 4435 13028 4459 13030
rect 4515 13028 4521 13030
rect 4213 13008 4521 13028
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3528 7886 3556 8434
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 3160 6322 3188 6802
rect 3252 6730 3280 7346
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2582 6012 2890 6032
rect 2582 6010 2588 6012
rect 2644 6010 2668 6012
rect 2724 6010 2748 6012
rect 2804 6010 2828 6012
rect 2884 6010 2890 6012
rect 2644 5958 2646 6010
rect 2826 5958 2828 6010
rect 2582 5956 2588 5958
rect 2644 5956 2668 5958
rect 2724 5956 2748 5958
rect 2804 5956 2828 5958
rect 2884 5956 2890 5958
rect 2582 5936 2890 5956
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2608 5012 2636 5238
rect 2872 5228 2924 5234
rect 2976 5216 3004 6190
rect 2924 5188 3004 5216
rect 3056 5228 3108 5234
rect 2872 5170 2924 5176
rect 3056 5170 3108 5176
rect 2884 5012 2912 5170
rect 2516 4984 2912 5012
rect 2964 5024 3016 5030
rect 2516 4622 2544 4984
rect 2964 4966 3016 4972
rect 2582 4924 2890 4944
rect 2582 4922 2588 4924
rect 2644 4922 2668 4924
rect 2724 4922 2748 4924
rect 2804 4922 2828 4924
rect 2884 4922 2890 4924
rect 2644 4870 2646 4922
rect 2826 4870 2828 4922
rect 2582 4868 2588 4870
rect 2644 4868 2668 4870
rect 2724 4868 2748 4870
rect 2804 4868 2828 4870
rect 2884 4868 2890 4870
rect 2582 4848 2890 4868
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2884 4078 2912 4422
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2332 3641 2360 3878
rect 2582 3836 2890 3856
rect 2582 3834 2588 3836
rect 2644 3834 2668 3836
rect 2724 3834 2748 3836
rect 2804 3834 2828 3836
rect 2884 3834 2890 3836
rect 2644 3782 2646 3834
rect 2826 3782 2828 3834
rect 2582 3780 2588 3782
rect 2644 3780 2668 3782
rect 2724 3780 2748 3782
rect 2804 3780 2828 3782
rect 2884 3780 2890 3782
rect 2582 3760 2890 3780
rect 2318 3632 2374 3641
rect 2318 3567 2374 3576
rect 2976 3058 3004 4966
rect 3068 4826 3096 5170
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3160 2774 3188 5034
rect 3344 4758 3372 7142
rect 3988 6798 4016 12582
rect 4213 11996 4521 12016
rect 4213 11994 4219 11996
rect 4275 11994 4299 11996
rect 4355 11994 4379 11996
rect 4435 11994 4459 11996
rect 4515 11994 4521 11996
rect 4275 11942 4277 11994
rect 4457 11942 4459 11994
rect 4213 11940 4219 11942
rect 4275 11940 4299 11942
rect 4355 11940 4379 11942
rect 4435 11940 4459 11942
rect 4515 11940 4521 11942
rect 4213 11920 4521 11940
rect 4213 10908 4521 10928
rect 4213 10906 4219 10908
rect 4275 10906 4299 10908
rect 4355 10906 4379 10908
rect 4435 10906 4459 10908
rect 4515 10906 4521 10908
rect 4275 10854 4277 10906
rect 4457 10854 4459 10906
rect 4213 10852 4219 10854
rect 4275 10852 4299 10854
rect 4355 10852 4379 10854
rect 4435 10852 4459 10854
rect 4515 10852 4521 10854
rect 4213 10832 4521 10852
rect 4213 9820 4521 9840
rect 4213 9818 4219 9820
rect 4275 9818 4299 9820
rect 4355 9818 4379 9820
rect 4435 9818 4459 9820
rect 4515 9818 4521 9820
rect 4275 9766 4277 9818
rect 4457 9766 4459 9818
rect 4213 9764 4219 9766
rect 4275 9764 4299 9766
rect 4355 9764 4379 9766
rect 4435 9764 4459 9766
rect 4515 9764 4521 9766
rect 4213 9744 4521 9764
rect 4213 8732 4521 8752
rect 4213 8730 4219 8732
rect 4275 8730 4299 8732
rect 4355 8730 4379 8732
rect 4435 8730 4459 8732
rect 4515 8730 4521 8732
rect 4275 8678 4277 8730
rect 4457 8678 4459 8730
rect 4213 8676 4219 8678
rect 4275 8676 4299 8678
rect 4355 8676 4379 8678
rect 4435 8676 4459 8678
rect 4515 8676 4521 8678
rect 4213 8656 4521 8676
rect 4213 7644 4521 7664
rect 4213 7642 4219 7644
rect 4275 7642 4299 7644
rect 4355 7642 4379 7644
rect 4435 7642 4459 7644
rect 4515 7642 4521 7644
rect 4275 7590 4277 7642
rect 4457 7590 4459 7642
rect 4213 7588 4219 7590
rect 4275 7588 4299 7590
rect 4355 7588 4379 7590
rect 4435 7588 4459 7590
rect 4515 7588 4521 7590
rect 4213 7568 4521 7588
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 5370 3924 6598
rect 4213 6556 4521 6576
rect 4213 6554 4219 6556
rect 4275 6554 4299 6556
rect 4355 6554 4379 6556
rect 4435 6554 4459 6556
rect 4515 6554 4521 6556
rect 4275 6502 4277 6554
rect 4457 6502 4459 6554
rect 4213 6500 4219 6502
rect 4275 6500 4299 6502
rect 4355 6500 4379 6502
rect 4435 6500 4459 6502
rect 4515 6500 4521 6502
rect 4213 6480 4521 6500
rect 4632 5914 4660 27950
rect 4724 5914 4752 28494
rect 4816 7886 4844 34886
rect 4908 23186 4936 50866
rect 4988 49768 5040 49774
rect 4988 49710 5040 49716
rect 5000 37194 5028 49710
rect 5172 40656 5224 40662
rect 5172 40598 5224 40604
rect 5080 40588 5132 40594
rect 5080 40530 5132 40536
rect 5092 39953 5120 40530
rect 5078 39944 5134 39953
rect 5078 39879 5134 39888
rect 5080 39840 5132 39846
rect 5080 39782 5132 39788
rect 5092 38962 5120 39782
rect 5080 38956 5132 38962
rect 5080 38898 5132 38904
rect 4988 37188 5040 37194
rect 4988 37130 5040 37136
rect 4988 36236 5040 36242
rect 4988 36178 5040 36184
rect 5000 34746 5028 36178
rect 5092 35578 5120 38898
rect 5184 36038 5212 40598
rect 5276 39574 5304 51046
rect 5368 40594 5396 65078
rect 5540 55208 5592 55214
rect 5540 55150 5592 55156
rect 5448 52420 5500 52426
rect 5448 52362 5500 52368
rect 5460 49706 5488 52362
rect 5448 49700 5500 49706
rect 5448 49642 5500 49648
rect 5356 40588 5408 40594
rect 5356 40530 5408 40536
rect 5356 40180 5408 40186
rect 5356 40122 5408 40128
rect 5264 39568 5316 39574
rect 5264 39510 5316 39516
rect 5262 39400 5318 39409
rect 5262 39335 5318 39344
rect 5172 36032 5224 36038
rect 5172 35974 5224 35980
rect 5276 35834 5304 39335
rect 5368 35873 5396 40122
rect 5354 35864 5410 35873
rect 5264 35828 5316 35834
rect 5354 35799 5410 35808
rect 5264 35770 5316 35776
rect 5460 35714 5488 49642
rect 5552 39914 5580 55150
rect 5540 39908 5592 39914
rect 5540 39850 5592 39856
rect 5644 38536 5672 74258
rect 5845 73468 6153 73488
rect 5845 73466 5851 73468
rect 5907 73466 5931 73468
rect 5987 73466 6011 73468
rect 6067 73466 6091 73468
rect 6147 73466 6153 73468
rect 5907 73414 5909 73466
rect 6089 73414 6091 73466
rect 5845 73412 5851 73414
rect 5907 73412 5931 73414
rect 5987 73412 6011 73414
rect 6067 73412 6091 73414
rect 6147 73412 6153 73414
rect 5845 73392 6153 73412
rect 5724 72480 5776 72486
rect 5724 72422 5776 72428
rect 5368 35686 5488 35714
rect 5552 38508 5672 38536
rect 5092 35550 5304 35578
rect 5172 35488 5224 35494
rect 5078 35456 5134 35465
rect 5172 35430 5224 35436
rect 5078 35391 5134 35400
rect 4988 34740 5040 34746
rect 4988 34682 5040 34688
rect 4988 34536 5040 34542
rect 4988 34478 5040 34484
rect 4896 23180 4948 23186
rect 4896 23122 4948 23128
rect 5000 8498 5028 34478
rect 5092 28218 5120 35391
rect 5184 30326 5212 35430
rect 5172 30320 5224 30326
rect 5172 30262 5224 30268
rect 5172 30048 5224 30054
rect 5172 29990 5224 29996
rect 5080 28212 5132 28218
rect 5080 28154 5132 28160
rect 5184 11082 5212 29990
rect 5276 17338 5304 35550
rect 5368 35494 5396 35686
rect 5448 35624 5500 35630
rect 5448 35566 5500 35572
rect 5356 35488 5408 35494
rect 5356 35430 5408 35436
rect 5356 34740 5408 34746
rect 5356 34682 5408 34688
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5368 8430 5396 34682
rect 5460 30938 5488 35566
rect 5552 35562 5580 38508
rect 5632 38208 5684 38214
rect 5632 38150 5684 38156
rect 5540 35556 5592 35562
rect 5540 35498 5592 35504
rect 5540 31952 5592 31958
rect 5540 31894 5592 31900
rect 5448 30932 5500 30938
rect 5448 30874 5500 30880
rect 5448 30592 5500 30598
rect 5448 30534 5500 30540
rect 5460 12646 5488 30534
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5552 7954 5580 31894
rect 5644 14482 5672 38150
rect 5736 34202 5764 72422
rect 5845 72380 6153 72400
rect 5845 72378 5851 72380
rect 5907 72378 5931 72380
rect 5987 72378 6011 72380
rect 6067 72378 6091 72380
rect 6147 72378 6153 72380
rect 5907 72326 5909 72378
rect 6089 72326 6091 72378
rect 5845 72324 5851 72326
rect 5907 72324 5931 72326
rect 5987 72324 6011 72326
rect 6067 72324 6091 72326
rect 6147 72324 6153 72326
rect 5845 72304 6153 72324
rect 6460 72004 6512 72010
rect 6460 71946 6512 71952
rect 5845 71292 6153 71312
rect 5845 71290 5851 71292
rect 5907 71290 5931 71292
rect 5987 71290 6011 71292
rect 6067 71290 6091 71292
rect 6147 71290 6153 71292
rect 5907 71238 5909 71290
rect 6089 71238 6091 71290
rect 5845 71236 5851 71238
rect 5907 71236 5931 71238
rect 5987 71236 6011 71238
rect 6067 71236 6091 71238
rect 6147 71236 6153 71238
rect 5845 71216 6153 71236
rect 5845 70204 6153 70224
rect 5845 70202 5851 70204
rect 5907 70202 5931 70204
rect 5987 70202 6011 70204
rect 6067 70202 6091 70204
rect 6147 70202 6153 70204
rect 5907 70150 5909 70202
rect 6089 70150 6091 70202
rect 5845 70148 5851 70150
rect 5907 70148 5931 70150
rect 5987 70148 6011 70150
rect 6067 70148 6091 70150
rect 6147 70148 6153 70150
rect 5845 70128 6153 70148
rect 5845 69116 6153 69136
rect 5845 69114 5851 69116
rect 5907 69114 5931 69116
rect 5987 69114 6011 69116
rect 6067 69114 6091 69116
rect 6147 69114 6153 69116
rect 5907 69062 5909 69114
rect 6089 69062 6091 69114
rect 5845 69060 5851 69062
rect 5907 69060 5931 69062
rect 5987 69060 6011 69062
rect 6067 69060 6091 69062
rect 6147 69060 6153 69062
rect 5845 69040 6153 69060
rect 6184 69012 6236 69018
rect 6184 68954 6236 68960
rect 5845 68028 6153 68048
rect 5845 68026 5851 68028
rect 5907 68026 5931 68028
rect 5987 68026 6011 68028
rect 6067 68026 6091 68028
rect 6147 68026 6153 68028
rect 5907 67974 5909 68026
rect 6089 67974 6091 68026
rect 5845 67972 5851 67974
rect 5907 67972 5931 67974
rect 5987 67972 6011 67974
rect 6067 67972 6091 67974
rect 6147 67972 6153 67974
rect 5845 67952 6153 67972
rect 5845 66940 6153 66960
rect 5845 66938 5851 66940
rect 5907 66938 5931 66940
rect 5987 66938 6011 66940
rect 6067 66938 6091 66940
rect 6147 66938 6153 66940
rect 5907 66886 5909 66938
rect 6089 66886 6091 66938
rect 5845 66884 5851 66886
rect 5907 66884 5931 66886
rect 5987 66884 6011 66886
rect 6067 66884 6091 66886
rect 6147 66884 6153 66886
rect 5845 66864 6153 66884
rect 5845 65852 6153 65872
rect 5845 65850 5851 65852
rect 5907 65850 5931 65852
rect 5987 65850 6011 65852
rect 6067 65850 6091 65852
rect 6147 65850 6153 65852
rect 5907 65798 5909 65850
rect 6089 65798 6091 65850
rect 5845 65796 5851 65798
rect 5907 65796 5931 65798
rect 5987 65796 6011 65798
rect 6067 65796 6091 65798
rect 6147 65796 6153 65798
rect 5845 65776 6153 65796
rect 5845 64764 6153 64784
rect 5845 64762 5851 64764
rect 5907 64762 5931 64764
rect 5987 64762 6011 64764
rect 6067 64762 6091 64764
rect 6147 64762 6153 64764
rect 5907 64710 5909 64762
rect 6089 64710 6091 64762
rect 5845 64708 5851 64710
rect 5907 64708 5931 64710
rect 5987 64708 6011 64710
rect 6067 64708 6091 64710
rect 6147 64708 6153 64710
rect 5845 64688 6153 64708
rect 5845 63676 6153 63696
rect 5845 63674 5851 63676
rect 5907 63674 5931 63676
rect 5987 63674 6011 63676
rect 6067 63674 6091 63676
rect 6147 63674 6153 63676
rect 5907 63622 5909 63674
rect 6089 63622 6091 63674
rect 5845 63620 5851 63622
rect 5907 63620 5931 63622
rect 5987 63620 6011 63622
rect 6067 63620 6091 63622
rect 6147 63620 6153 63622
rect 5845 63600 6153 63620
rect 5845 62588 6153 62608
rect 5845 62586 5851 62588
rect 5907 62586 5931 62588
rect 5987 62586 6011 62588
rect 6067 62586 6091 62588
rect 6147 62586 6153 62588
rect 5907 62534 5909 62586
rect 6089 62534 6091 62586
rect 5845 62532 5851 62534
rect 5907 62532 5931 62534
rect 5987 62532 6011 62534
rect 6067 62532 6091 62534
rect 6147 62532 6153 62534
rect 5845 62512 6153 62532
rect 5845 61500 6153 61520
rect 5845 61498 5851 61500
rect 5907 61498 5931 61500
rect 5987 61498 6011 61500
rect 6067 61498 6091 61500
rect 6147 61498 6153 61500
rect 5907 61446 5909 61498
rect 6089 61446 6091 61498
rect 5845 61444 5851 61446
rect 5907 61444 5931 61446
rect 5987 61444 6011 61446
rect 6067 61444 6091 61446
rect 6147 61444 6153 61446
rect 5845 61424 6153 61444
rect 5845 60412 6153 60432
rect 5845 60410 5851 60412
rect 5907 60410 5931 60412
rect 5987 60410 6011 60412
rect 6067 60410 6091 60412
rect 6147 60410 6153 60412
rect 5907 60358 5909 60410
rect 6089 60358 6091 60410
rect 5845 60356 5851 60358
rect 5907 60356 5931 60358
rect 5987 60356 6011 60358
rect 6067 60356 6091 60358
rect 6147 60356 6153 60358
rect 5845 60336 6153 60356
rect 5845 59324 6153 59344
rect 5845 59322 5851 59324
rect 5907 59322 5931 59324
rect 5987 59322 6011 59324
rect 6067 59322 6091 59324
rect 6147 59322 6153 59324
rect 5907 59270 5909 59322
rect 6089 59270 6091 59322
rect 5845 59268 5851 59270
rect 5907 59268 5931 59270
rect 5987 59268 6011 59270
rect 6067 59268 6091 59270
rect 6147 59268 6153 59270
rect 5845 59248 6153 59268
rect 5845 58236 6153 58256
rect 5845 58234 5851 58236
rect 5907 58234 5931 58236
rect 5987 58234 6011 58236
rect 6067 58234 6091 58236
rect 6147 58234 6153 58236
rect 5907 58182 5909 58234
rect 6089 58182 6091 58234
rect 5845 58180 5851 58182
rect 5907 58180 5931 58182
rect 5987 58180 6011 58182
rect 6067 58180 6091 58182
rect 6147 58180 6153 58182
rect 5845 58160 6153 58180
rect 5845 57148 6153 57168
rect 5845 57146 5851 57148
rect 5907 57146 5931 57148
rect 5987 57146 6011 57148
rect 6067 57146 6091 57148
rect 6147 57146 6153 57148
rect 5907 57094 5909 57146
rect 6089 57094 6091 57146
rect 5845 57092 5851 57094
rect 5907 57092 5931 57094
rect 5987 57092 6011 57094
rect 6067 57092 6091 57094
rect 6147 57092 6153 57094
rect 5845 57072 6153 57092
rect 5816 56432 5868 56438
rect 5816 56374 5868 56380
rect 5828 56273 5856 56374
rect 5814 56264 5870 56273
rect 5814 56199 5870 56208
rect 5845 56060 6153 56080
rect 5845 56058 5851 56060
rect 5907 56058 5931 56060
rect 5987 56058 6011 56060
rect 6067 56058 6091 56060
rect 6147 56058 6153 56060
rect 5907 56006 5909 56058
rect 6089 56006 6091 56058
rect 5845 56004 5851 56006
rect 5907 56004 5931 56006
rect 5987 56004 6011 56006
rect 6067 56004 6091 56006
rect 6147 56004 6153 56006
rect 5845 55984 6153 56004
rect 5845 54972 6153 54992
rect 5845 54970 5851 54972
rect 5907 54970 5931 54972
rect 5987 54970 6011 54972
rect 6067 54970 6091 54972
rect 6147 54970 6153 54972
rect 5907 54918 5909 54970
rect 6089 54918 6091 54970
rect 5845 54916 5851 54918
rect 5907 54916 5931 54918
rect 5987 54916 6011 54918
rect 6067 54916 6091 54918
rect 6147 54916 6153 54918
rect 5845 54896 6153 54916
rect 5845 53884 6153 53904
rect 5845 53882 5851 53884
rect 5907 53882 5931 53884
rect 5987 53882 6011 53884
rect 6067 53882 6091 53884
rect 6147 53882 6153 53884
rect 5907 53830 5909 53882
rect 6089 53830 6091 53882
rect 5845 53828 5851 53830
rect 5907 53828 5931 53830
rect 5987 53828 6011 53830
rect 6067 53828 6091 53830
rect 6147 53828 6153 53830
rect 5845 53808 6153 53828
rect 5845 52796 6153 52816
rect 5845 52794 5851 52796
rect 5907 52794 5931 52796
rect 5987 52794 6011 52796
rect 6067 52794 6091 52796
rect 6147 52794 6153 52796
rect 5907 52742 5909 52794
rect 6089 52742 6091 52794
rect 5845 52740 5851 52742
rect 5907 52740 5931 52742
rect 5987 52740 6011 52742
rect 6067 52740 6091 52742
rect 6147 52740 6153 52742
rect 5845 52720 6153 52740
rect 5845 51708 6153 51728
rect 5845 51706 5851 51708
rect 5907 51706 5931 51708
rect 5987 51706 6011 51708
rect 6067 51706 6091 51708
rect 6147 51706 6153 51708
rect 5907 51654 5909 51706
rect 6089 51654 6091 51706
rect 5845 51652 5851 51654
rect 5907 51652 5931 51654
rect 5987 51652 6011 51654
rect 6067 51652 6091 51654
rect 6147 51652 6153 51654
rect 5845 51632 6153 51652
rect 5816 51468 5868 51474
rect 5816 51410 5868 51416
rect 5828 51377 5856 51410
rect 5814 51368 5870 51377
rect 5814 51303 5870 51312
rect 5845 50620 6153 50640
rect 5845 50618 5851 50620
rect 5907 50618 5931 50620
rect 5987 50618 6011 50620
rect 6067 50618 6091 50620
rect 6147 50618 6153 50620
rect 5907 50566 5909 50618
rect 6089 50566 6091 50618
rect 5845 50564 5851 50566
rect 5907 50564 5931 50566
rect 5987 50564 6011 50566
rect 6067 50564 6091 50566
rect 6147 50564 6153 50566
rect 5845 50544 6153 50564
rect 5845 49532 6153 49552
rect 5845 49530 5851 49532
rect 5907 49530 5931 49532
rect 5987 49530 6011 49532
rect 6067 49530 6091 49532
rect 6147 49530 6153 49532
rect 5907 49478 5909 49530
rect 6089 49478 6091 49530
rect 5845 49476 5851 49478
rect 5907 49476 5931 49478
rect 5987 49476 6011 49478
rect 6067 49476 6091 49478
rect 6147 49476 6153 49478
rect 5845 49456 6153 49476
rect 5845 48444 6153 48464
rect 5845 48442 5851 48444
rect 5907 48442 5931 48444
rect 5987 48442 6011 48444
rect 6067 48442 6091 48444
rect 6147 48442 6153 48444
rect 5907 48390 5909 48442
rect 6089 48390 6091 48442
rect 5845 48388 5851 48390
rect 5907 48388 5931 48390
rect 5987 48388 6011 48390
rect 6067 48388 6091 48390
rect 6147 48388 6153 48390
rect 5845 48368 6153 48388
rect 5845 47356 6153 47376
rect 5845 47354 5851 47356
rect 5907 47354 5931 47356
rect 5987 47354 6011 47356
rect 6067 47354 6091 47356
rect 6147 47354 6153 47356
rect 5907 47302 5909 47354
rect 6089 47302 6091 47354
rect 5845 47300 5851 47302
rect 5907 47300 5931 47302
rect 5987 47300 6011 47302
rect 6067 47300 6091 47302
rect 6147 47300 6153 47302
rect 5845 47280 6153 47300
rect 5845 46268 6153 46288
rect 5845 46266 5851 46268
rect 5907 46266 5931 46268
rect 5987 46266 6011 46268
rect 6067 46266 6091 46268
rect 6147 46266 6153 46268
rect 5907 46214 5909 46266
rect 6089 46214 6091 46266
rect 5845 46212 5851 46214
rect 5907 46212 5931 46214
rect 5987 46212 6011 46214
rect 6067 46212 6091 46214
rect 6147 46212 6153 46214
rect 5845 46192 6153 46212
rect 5845 45180 6153 45200
rect 5845 45178 5851 45180
rect 5907 45178 5931 45180
rect 5987 45178 6011 45180
rect 6067 45178 6091 45180
rect 6147 45178 6153 45180
rect 5907 45126 5909 45178
rect 6089 45126 6091 45178
rect 5845 45124 5851 45126
rect 5907 45124 5931 45126
rect 5987 45124 6011 45126
rect 6067 45124 6091 45126
rect 6147 45124 6153 45126
rect 5845 45104 6153 45124
rect 5845 44092 6153 44112
rect 5845 44090 5851 44092
rect 5907 44090 5931 44092
rect 5987 44090 6011 44092
rect 6067 44090 6091 44092
rect 6147 44090 6153 44092
rect 5907 44038 5909 44090
rect 6089 44038 6091 44090
rect 5845 44036 5851 44038
rect 5907 44036 5931 44038
rect 5987 44036 6011 44038
rect 6067 44036 6091 44038
rect 6147 44036 6153 44038
rect 5845 44016 6153 44036
rect 5845 43004 6153 43024
rect 5845 43002 5851 43004
rect 5907 43002 5931 43004
rect 5987 43002 6011 43004
rect 6067 43002 6091 43004
rect 6147 43002 6153 43004
rect 5907 42950 5909 43002
rect 6089 42950 6091 43002
rect 5845 42948 5851 42950
rect 5907 42948 5931 42950
rect 5987 42948 6011 42950
rect 6067 42948 6091 42950
rect 6147 42948 6153 42950
rect 5845 42928 6153 42948
rect 5845 41916 6153 41936
rect 5845 41914 5851 41916
rect 5907 41914 5931 41916
rect 5987 41914 6011 41916
rect 6067 41914 6091 41916
rect 6147 41914 6153 41916
rect 5907 41862 5909 41914
rect 6089 41862 6091 41914
rect 5845 41860 5851 41862
rect 5907 41860 5931 41862
rect 5987 41860 6011 41862
rect 6067 41860 6091 41862
rect 6147 41860 6153 41862
rect 5845 41840 6153 41860
rect 5845 40828 6153 40848
rect 5845 40826 5851 40828
rect 5907 40826 5931 40828
rect 5987 40826 6011 40828
rect 6067 40826 6091 40828
rect 6147 40826 6153 40828
rect 5907 40774 5909 40826
rect 6089 40774 6091 40826
rect 5845 40772 5851 40774
rect 5907 40772 5931 40774
rect 5987 40772 6011 40774
rect 6067 40772 6091 40774
rect 6147 40772 6153 40774
rect 5845 40752 6153 40772
rect 5845 39740 6153 39760
rect 5845 39738 5851 39740
rect 5907 39738 5931 39740
rect 5987 39738 6011 39740
rect 6067 39738 6091 39740
rect 6147 39738 6153 39740
rect 5907 39686 5909 39738
rect 6089 39686 6091 39738
rect 5845 39684 5851 39686
rect 5907 39684 5931 39686
rect 5987 39684 6011 39686
rect 6067 39684 6091 39686
rect 6147 39684 6153 39686
rect 5845 39664 6153 39684
rect 5845 38652 6153 38672
rect 5845 38650 5851 38652
rect 5907 38650 5931 38652
rect 5987 38650 6011 38652
rect 6067 38650 6091 38652
rect 6147 38650 6153 38652
rect 5907 38598 5909 38650
rect 6089 38598 6091 38650
rect 5845 38596 5851 38598
rect 5907 38596 5931 38598
rect 5987 38596 6011 38598
rect 6067 38596 6091 38598
rect 6147 38596 6153 38598
rect 5845 38576 6153 38596
rect 6196 38010 6224 68954
rect 6276 50176 6328 50182
rect 6276 50118 6328 50124
rect 6184 38004 6236 38010
rect 6184 37946 6236 37952
rect 6184 37664 6236 37670
rect 6184 37606 6236 37612
rect 5845 37564 6153 37584
rect 5845 37562 5851 37564
rect 5907 37562 5931 37564
rect 5987 37562 6011 37564
rect 6067 37562 6091 37564
rect 6147 37562 6153 37564
rect 5907 37510 5909 37562
rect 6089 37510 6091 37562
rect 5845 37508 5851 37510
rect 5907 37508 5931 37510
rect 5987 37508 6011 37510
rect 6067 37508 6091 37510
rect 6147 37508 6153 37510
rect 5845 37488 6153 37508
rect 5845 36476 6153 36496
rect 5845 36474 5851 36476
rect 5907 36474 5931 36476
rect 5987 36474 6011 36476
rect 6067 36474 6091 36476
rect 6147 36474 6153 36476
rect 5907 36422 5909 36474
rect 6089 36422 6091 36474
rect 5845 36420 5851 36422
rect 5907 36420 5931 36422
rect 5987 36420 6011 36422
rect 6067 36420 6091 36422
rect 6147 36420 6153 36422
rect 5845 36400 6153 36420
rect 5845 35388 6153 35408
rect 5845 35386 5851 35388
rect 5907 35386 5931 35388
rect 5987 35386 6011 35388
rect 6067 35386 6091 35388
rect 6147 35386 6153 35388
rect 5907 35334 5909 35386
rect 6089 35334 6091 35386
rect 5845 35332 5851 35334
rect 5907 35332 5931 35334
rect 5987 35332 6011 35334
rect 6067 35332 6091 35334
rect 6147 35332 6153 35334
rect 5845 35312 6153 35332
rect 5845 34300 6153 34320
rect 5845 34298 5851 34300
rect 5907 34298 5931 34300
rect 5987 34298 6011 34300
rect 6067 34298 6091 34300
rect 6147 34298 6153 34300
rect 5907 34246 5909 34298
rect 6089 34246 6091 34298
rect 5845 34244 5851 34246
rect 5907 34244 5931 34246
rect 5987 34244 6011 34246
rect 6067 34244 6091 34246
rect 6147 34244 6153 34246
rect 5845 34224 6153 34244
rect 5724 34196 5776 34202
rect 5724 34138 5776 34144
rect 5845 33212 6153 33232
rect 5845 33210 5851 33212
rect 5907 33210 5931 33212
rect 5987 33210 6011 33212
rect 6067 33210 6091 33212
rect 6147 33210 6153 33212
rect 5907 33158 5909 33210
rect 6089 33158 6091 33210
rect 5845 33156 5851 33158
rect 5907 33156 5931 33158
rect 5987 33156 6011 33158
rect 6067 33156 6091 33158
rect 6147 33156 6153 33158
rect 5845 33136 6153 33156
rect 5845 32124 6153 32144
rect 5845 32122 5851 32124
rect 5907 32122 5931 32124
rect 5987 32122 6011 32124
rect 6067 32122 6091 32124
rect 6147 32122 6153 32124
rect 5907 32070 5909 32122
rect 6089 32070 6091 32122
rect 5845 32068 5851 32070
rect 5907 32068 5931 32070
rect 5987 32068 6011 32070
rect 6067 32068 6091 32070
rect 6147 32068 6153 32070
rect 5845 32048 6153 32068
rect 5845 31036 6153 31056
rect 5845 31034 5851 31036
rect 5907 31034 5931 31036
rect 5987 31034 6011 31036
rect 6067 31034 6091 31036
rect 6147 31034 6153 31036
rect 5907 30982 5909 31034
rect 6089 30982 6091 31034
rect 5845 30980 5851 30982
rect 5907 30980 5931 30982
rect 5987 30980 6011 30982
rect 6067 30980 6091 30982
rect 6147 30980 6153 30982
rect 5845 30960 6153 30980
rect 5845 29948 6153 29968
rect 5845 29946 5851 29948
rect 5907 29946 5931 29948
rect 5987 29946 6011 29948
rect 6067 29946 6091 29948
rect 6147 29946 6153 29948
rect 5907 29894 5909 29946
rect 6089 29894 6091 29946
rect 5845 29892 5851 29894
rect 5907 29892 5931 29894
rect 5987 29892 6011 29894
rect 6067 29892 6091 29894
rect 6147 29892 6153 29894
rect 5845 29872 6153 29892
rect 5845 28860 6153 28880
rect 5845 28858 5851 28860
rect 5907 28858 5931 28860
rect 5987 28858 6011 28860
rect 6067 28858 6091 28860
rect 6147 28858 6153 28860
rect 5907 28806 5909 28858
rect 6089 28806 6091 28858
rect 5845 28804 5851 28806
rect 5907 28804 5931 28806
rect 5987 28804 6011 28806
rect 6067 28804 6091 28806
rect 6147 28804 6153 28806
rect 5845 28784 6153 28804
rect 5845 27772 6153 27792
rect 5845 27770 5851 27772
rect 5907 27770 5931 27772
rect 5987 27770 6011 27772
rect 6067 27770 6091 27772
rect 6147 27770 6153 27772
rect 5907 27718 5909 27770
rect 6089 27718 6091 27770
rect 5845 27716 5851 27718
rect 5907 27716 5931 27718
rect 5987 27716 6011 27718
rect 6067 27716 6091 27718
rect 6147 27716 6153 27718
rect 5845 27696 6153 27716
rect 5845 26684 6153 26704
rect 5845 26682 5851 26684
rect 5907 26682 5931 26684
rect 5987 26682 6011 26684
rect 6067 26682 6091 26684
rect 6147 26682 6153 26684
rect 5907 26630 5909 26682
rect 6089 26630 6091 26682
rect 5845 26628 5851 26630
rect 5907 26628 5931 26630
rect 5987 26628 6011 26630
rect 6067 26628 6091 26630
rect 6147 26628 6153 26630
rect 5845 26608 6153 26628
rect 5845 25596 6153 25616
rect 5845 25594 5851 25596
rect 5907 25594 5931 25596
rect 5987 25594 6011 25596
rect 6067 25594 6091 25596
rect 6147 25594 6153 25596
rect 5907 25542 5909 25594
rect 6089 25542 6091 25594
rect 5845 25540 5851 25542
rect 5907 25540 5931 25542
rect 5987 25540 6011 25542
rect 6067 25540 6091 25542
rect 6147 25540 6153 25542
rect 5845 25520 6153 25540
rect 5845 24508 6153 24528
rect 5845 24506 5851 24508
rect 5907 24506 5931 24508
rect 5987 24506 6011 24508
rect 6067 24506 6091 24508
rect 6147 24506 6153 24508
rect 5907 24454 5909 24506
rect 6089 24454 6091 24506
rect 5845 24452 5851 24454
rect 5907 24452 5931 24454
rect 5987 24452 6011 24454
rect 6067 24452 6091 24454
rect 6147 24452 6153 24454
rect 5845 24432 6153 24452
rect 5845 23420 6153 23440
rect 5845 23418 5851 23420
rect 5907 23418 5931 23420
rect 5987 23418 6011 23420
rect 6067 23418 6091 23420
rect 6147 23418 6153 23420
rect 5907 23366 5909 23418
rect 6089 23366 6091 23418
rect 5845 23364 5851 23366
rect 5907 23364 5931 23366
rect 5987 23364 6011 23366
rect 6067 23364 6091 23366
rect 6147 23364 6153 23366
rect 5845 23344 6153 23364
rect 5845 22332 6153 22352
rect 5845 22330 5851 22332
rect 5907 22330 5931 22332
rect 5987 22330 6011 22332
rect 6067 22330 6091 22332
rect 6147 22330 6153 22332
rect 5907 22278 5909 22330
rect 6089 22278 6091 22330
rect 5845 22276 5851 22278
rect 5907 22276 5931 22278
rect 5987 22276 6011 22278
rect 6067 22276 6091 22278
rect 6147 22276 6153 22278
rect 5845 22256 6153 22276
rect 5845 21244 6153 21264
rect 5845 21242 5851 21244
rect 5907 21242 5931 21244
rect 5987 21242 6011 21244
rect 6067 21242 6091 21244
rect 6147 21242 6153 21244
rect 5907 21190 5909 21242
rect 6089 21190 6091 21242
rect 5845 21188 5851 21190
rect 5907 21188 5931 21190
rect 5987 21188 6011 21190
rect 6067 21188 6091 21190
rect 6147 21188 6153 21190
rect 5845 21168 6153 21188
rect 5845 20156 6153 20176
rect 5845 20154 5851 20156
rect 5907 20154 5931 20156
rect 5987 20154 6011 20156
rect 6067 20154 6091 20156
rect 6147 20154 6153 20156
rect 5907 20102 5909 20154
rect 6089 20102 6091 20154
rect 5845 20100 5851 20102
rect 5907 20100 5931 20102
rect 5987 20100 6011 20102
rect 6067 20100 6091 20102
rect 6147 20100 6153 20102
rect 5845 20080 6153 20100
rect 5845 19068 6153 19088
rect 5845 19066 5851 19068
rect 5907 19066 5931 19068
rect 5987 19066 6011 19068
rect 6067 19066 6091 19068
rect 6147 19066 6153 19068
rect 5907 19014 5909 19066
rect 6089 19014 6091 19066
rect 5845 19012 5851 19014
rect 5907 19012 5931 19014
rect 5987 19012 6011 19014
rect 6067 19012 6091 19014
rect 6147 19012 6153 19014
rect 5845 18992 6153 19012
rect 5845 17980 6153 18000
rect 5845 17978 5851 17980
rect 5907 17978 5931 17980
rect 5987 17978 6011 17980
rect 6067 17978 6091 17980
rect 6147 17978 6153 17980
rect 5907 17926 5909 17978
rect 6089 17926 6091 17978
rect 5845 17924 5851 17926
rect 5907 17924 5931 17926
rect 5987 17924 6011 17926
rect 6067 17924 6091 17926
rect 6147 17924 6153 17926
rect 5845 17904 6153 17924
rect 5845 16892 6153 16912
rect 5845 16890 5851 16892
rect 5907 16890 5931 16892
rect 5987 16890 6011 16892
rect 6067 16890 6091 16892
rect 6147 16890 6153 16892
rect 5907 16838 5909 16890
rect 6089 16838 6091 16890
rect 5845 16836 5851 16838
rect 5907 16836 5931 16838
rect 5987 16836 6011 16838
rect 6067 16836 6091 16838
rect 6147 16836 6153 16838
rect 5845 16816 6153 16836
rect 5845 15804 6153 15824
rect 5845 15802 5851 15804
rect 5907 15802 5931 15804
rect 5987 15802 6011 15804
rect 6067 15802 6091 15804
rect 6147 15802 6153 15804
rect 5907 15750 5909 15802
rect 6089 15750 6091 15802
rect 5845 15748 5851 15750
rect 5907 15748 5931 15750
rect 5987 15748 6011 15750
rect 6067 15748 6091 15750
rect 6147 15748 6153 15750
rect 5845 15728 6153 15748
rect 6196 14958 6224 37606
rect 6288 24206 6316 50118
rect 6368 44804 6420 44810
rect 6368 44746 6420 44752
rect 6276 24200 6328 24206
rect 6276 24142 6328 24148
rect 6380 17202 6408 44746
rect 6472 41206 6500 71946
rect 6460 41200 6512 41206
rect 6460 41142 6512 41148
rect 6564 41018 6592 74870
rect 7477 74012 7785 74032
rect 7477 74010 7483 74012
rect 7539 74010 7563 74012
rect 7619 74010 7643 74012
rect 7699 74010 7723 74012
rect 7779 74010 7785 74012
rect 7539 73958 7541 74010
rect 7721 73958 7723 74010
rect 7477 73956 7483 73958
rect 7539 73956 7563 73958
rect 7619 73956 7643 73958
rect 7699 73956 7723 73958
rect 7779 73956 7785 73958
rect 7477 73936 7785 73956
rect 8312 73914 8340 76978
rect 9109 76732 9417 76752
rect 9109 76730 9115 76732
rect 9171 76730 9195 76732
rect 9251 76730 9275 76732
rect 9331 76730 9355 76732
rect 9411 76730 9417 76732
rect 9171 76678 9173 76730
rect 9353 76678 9355 76730
rect 9109 76676 9115 76678
rect 9171 76676 9195 76678
rect 9251 76676 9275 76678
rect 9331 76676 9355 76678
rect 9411 76676 9417 76678
rect 9109 76656 9417 76676
rect 9109 75644 9417 75664
rect 9109 75642 9115 75644
rect 9171 75642 9195 75644
rect 9251 75642 9275 75644
rect 9331 75642 9355 75644
rect 9411 75642 9417 75644
rect 9171 75590 9173 75642
rect 9353 75590 9355 75642
rect 9109 75588 9115 75590
rect 9171 75588 9195 75590
rect 9251 75588 9275 75590
rect 9331 75588 9355 75590
rect 9411 75588 9417 75590
rect 9109 75568 9417 75588
rect 9109 74556 9417 74576
rect 9109 74554 9115 74556
rect 9171 74554 9195 74556
rect 9251 74554 9275 74556
rect 9331 74554 9355 74556
rect 9411 74554 9417 74556
rect 9171 74502 9173 74554
rect 9353 74502 9355 74554
rect 9109 74500 9115 74502
rect 9171 74500 9195 74502
rect 9251 74500 9275 74502
rect 9331 74500 9355 74502
rect 9411 74500 9417 74502
rect 9109 74480 9417 74500
rect 9692 74390 9720 76978
rect 10048 76832 10100 76838
rect 10048 76774 10100 76780
rect 10060 76537 10088 76774
rect 10046 76528 10102 76537
rect 10046 76463 10102 76472
rect 9772 76424 9824 76430
rect 9772 76366 9824 76372
rect 9680 74384 9732 74390
rect 9680 74326 9732 74332
rect 8300 73908 8352 73914
rect 8300 73850 8352 73856
rect 9784 73846 9812 76366
rect 10048 75744 10100 75750
rect 10046 75712 10048 75721
rect 10100 75712 10102 75721
rect 10046 75647 10102 75656
rect 9864 75336 9916 75342
rect 9864 75278 9916 75284
rect 9876 74458 9904 75278
rect 10048 75200 10100 75206
rect 10048 75142 10100 75148
rect 10060 75041 10088 75142
rect 10046 75032 10102 75041
rect 10046 74967 10102 74976
rect 9864 74452 9916 74458
rect 9864 74394 9916 74400
rect 9864 74248 9916 74254
rect 9864 74190 9916 74196
rect 10046 74216 10102 74225
rect 9772 73840 9824 73846
rect 9772 73782 9824 73788
rect 9876 73574 9904 74190
rect 10046 74151 10102 74160
rect 10060 74118 10088 74151
rect 10048 74112 10100 74118
rect 10048 74054 10100 74060
rect 9864 73568 9916 73574
rect 10048 73568 10100 73574
rect 9864 73510 9916 73516
rect 10046 73536 10048 73545
rect 10100 73536 10102 73545
rect 9109 73468 9417 73488
rect 10046 73471 10102 73480
rect 9109 73466 9115 73468
rect 9171 73466 9195 73468
rect 9251 73466 9275 73468
rect 9331 73466 9355 73468
rect 9411 73466 9417 73468
rect 9171 73414 9173 73466
rect 9353 73414 9355 73466
rect 9109 73412 9115 73414
rect 9171 73412 9195 73414
rect 9251 73412 9275 73414
rect 9331 73412 9355 73414
rect 9411 73412 9417 73414
rect 9109 73392 9417 73412
rect 10048 73024 10100 73030
rect 10048 72966 10100 72972
rect 7477 72924 7785 72944
rect 7477 72922 7483 72924
rect 7539 72922 7563 72924
rect 7619 72922 7643 72924
rect 7699 72922 7723 72924
rect 7779 72922 7785 72924
rect 7539 72870 7541 72922
rect 7721 72870 7723 72922
rect 7477 72868 7483 72870
rect 7539 72868 7563 72870
rect 7619 72868 7643 72870
rect 7699 72868 7723 72870
rect 7779 72868 7785 72870
rect 7477 72848 7785 72868
rect 10060 72729 10088 72966
rect 10046 72720 10102 72729
rect 10046 72655 10102 72664
rect 7012 72548 7064 72554
rect 7012 72490 7064 72496
rect 6644 65000 6696 65006
rect 6644 64942 6696 64948
rect 6656 41313 6684 64942
rect 6920 63300 6972 63306
rect 6920 63242 6972 63248
rect 6736 45280 6788 45286
rect 6736 45222 6788 45228
rect 6642 41304 6698 41313
rect 6642 41239 6698 41248
rect 6644 41200 6696 41206
rect 6644 41142 6696 41148
rect 6472 40990 6592 41018
rect 6472 37126 6500 40990
rect 6552 40928 6604 40934
rect 6552 40870 6604 40876
rect 6460 37120 6512 37126
rect 6460 37062 6512 37068
rect 6458 36952 6514 36961
rect 6458 36887 6514 36896
rect 6472 32298 6500 36887
rect 6460 32292 6512 32298
rect 6460 32234 6512 32240
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6564 16182 6592 40870
rect 6656 34678 6684 41142
rect 6644 34672 6696 34678
rect 6644 34614 6696 34620
rect 6748 18086 6776 45222
rect 6828 40384 6880 40390
rect 6828 40326 6880 40332
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6552 16176 6604 16182
rect 6552 16118 6604 16124
rect 6840 15502 6868 40326
rect 6932 31754 6960 63242
rect 7024 38486 7052 72490
rect 9109 72380 9417 72400
rect 9109 72378 9115 72380
rect 9171 72378 9195 72380
rect 9251 72378 9275 72380
rect 9331 72378 9355 72380
rect 9411 72378 9417 72380
rect 9171 72326 9173 72378
rect 9353 72326 9355 72378
rect 9109 72324 9115 72326
rect 9171 72324 9195 72326
rect 9251 72324 9275 72326
rect 9331 72324 9355 72326
rect 9411 72324 9417 72326
rect 9109 72304 9417 72324
rect 9864 71936 9916 71942
rect 10048 71936 10100 71942
rect 9864 71878 9916 71884
rect 10046 71904 10048 71913
rect 10100 71904 10102 71913
rect 7477 71836 7785 71856
rect 7477 71834 7483 71836
rect 7539 71834 7563 71836
rect 7619 71834 7643 71836
rect 7699 71834 7723 71836
rect 7779 71834 7785 71836
rect 7539 71782 7541 71834
rect 7721 71782 7723 71834
rect 7477 71780 7483 71782
rect 7539 71780 7563 71782
rect 7619 71780 7643 71782
rect 7699 71780 7723 71782
rect 7779 71780 7785 71782
rect 7477 71760 7785 71780
rect 9876 71602 9904 71878
rect 10046 71839 10102 71848
rect 9864 71596 9916 71602
rect 9864 71538 9916 71544
rect 9864 71392 9916 71398
rect 9864 71334 9916 71340
rect 10048 71392 10100 71398
rect 10048 71334 10100 71340
rect 9109 71292 9417 71312
rect 9109 71290 9115 71292
rect 9171 71290 9195 71292
rect 9251 71290 9275 71292
rect 9331 71290 9355 71292
rect 9411 71290 9417 71292
rect 9171 71238 9173 71290
rect 9353 71238 9355 71290
rect 9109 71236 9115 71238
rect 9171 71236 9195 71238
rect 9251 71236 9275 71238
rect 9331 71236 9355 71238
rect 9411 71236 9417 71238
rect 9109 71216 9417 71236
rect 7477 70748 7785 70768
rect 7477 70746 7483 70748
rect 7539 70746 7563 70748
rect 7619 70746 7643 70748
rect 7699 70746 7723 70748
rect 7779 70746 7785 70748
rect 7539 70694 7541 70746
rect 7721 70694 7723 70746
rect 7477 70692 7483 70694
rect 7539 70692 7563 70694
rect 7619 70692 7643 70694
rect 7699 70692 7723 70694
rect 7779 70692 7785 70694
rect 7477 70672 7785 70692
rect 9876 70514 9904 71334
rect 10060 71233 10088 71334
rect 10046 71224 10102 71233
rect 10046 71159 10102 71168
rect 10692 70644 10744 70650
rect 10692 70586 10744 70592
rect 9864 70508 9916 70514
rect 9864 70450 9916 70456
rect 10704 70417 10732 70586
rect 10690 70408 10746 70417
rect 10690 70343 10746 70352
rect 9109 70204 9417 70224
rect 9109 70202 9115 70204
rect 9171 70202 9195 70204
rect 9251 70202 9275 70204
rect 9331 70202 9355 70204
rect 9411 70202 9417 70204
rect 9171 70150 9173 70202
rect 9353 70150 9355 70202
rect 9109 70148 9115 70150
rect 9171 70148 9195 70150
rect 9251 70148 9275 70150
rect 9331 70148 9355 70150
rect 9411 70148 9417 70150
rect 9109 70128 9417 70148
rect 10048 69760 10100 69766
rect 10046 69728 10048 69737
rect 10100 69728 10102 69737
rect 7477 69660 7785 69680
rect 10046 69663 10102 69672
rect 7477 69658 7483 69660
rect 7539 69658 7563 69660
rect 7619 69658 7643 69660
rect 7699 69658 7723 69660
rect 7779 69658 7785 69660
rect 7539 69606 7541 69658
rect 7721 69606 7723 69658
rect 7477 69604 7483 69606
rect 7539 69604 7563 69606
rect 7619 69604 7643 69606
rect 7699 69604 7723 69606
rect 7779 69604 7785 69606
rect 7477 69584 7785 69604
rect 10048 69216 10100 69222
rect 10048 69158 10100 69164
rect 9109 69116 9417 69136
rect 9109 69114 9115 69116
rect 9171 69114 9195 69116
rect 9251 69114 9275 69116
rect 9331 69114 9355 69116
rect 9411 69114 9417 69116
rect 9171 69062 9173 69114
rect 9353 69062 9355 69114
rect 9109 69060 9115 69062
rect 9171 69060 9195 69062
rect 9251 69060 9275 69062
rect 9331 69060 9355 69062
rect 9411 69060 9417 69062
rect 9109 69040 9417 69060
rect 10060 68921 10088 69158
rect 10046 68912 10102 68921
rect 10046 68847 10102 68856
rect 7477 68572 7785 68592
rect 7477 68570 7483 68572
rect 7539 68570 7563 68572
rect 7619 68570 7643 68572
rect 7699 68570 7723 68572
rect 7779 68570 7785 68572
rect 7539 68518 7541 68570
rect 7721 68518 7723 68570
rect 7477 68516 7483 68518
rect 7539 68516 7563 68518
rect 7619 68516 7643 68518
rect 7699 68516 7723 68518
rect 7779 68516 7785 68518
rect 7477 68496 7785 68516
rect 9864 68332 9916 68338
rect 9864 68274 9916 68280
rect 9109 68028 9417 68048
rect 9109 68026 9115 68028
rect 9171 68026 9195 68028
rect 9251 68026 9275 68028
rect 9331 68026 9355 68028
rect 9411 68026 9417 68028
rect 9171 67974 9173 68026
rect 9353 67974 9355 68026
rect 9109 67972 9115 67974
rect 9171 67972 9195 67974
rect 9251 67972 9275 67974
rect 9331 67972 9355 67974
rect 9411 67972 9417 67974
rect 9109 67952 9417 67972
rect 9772 67720 9824 67726
rect 9772 67662 9824 67668
rect 7477 67484 7785 67504
rect 7477 67482 7483 67484
rect 7539 67482 7563 67484
rect 7619 67482 7643 67484
rect 7699 67482 7723 67484
rect 7779 67482 7785 67484
rect 7539 67430 7541 67482
rect 7721 67430 7723 67482
rect 7477 67428 7483 67430
rect 7539 67428 7563 67430
rect 7619 67428 7643 67430
rect 7699 67428 7723 67430
rect 7779 67428 7785 67430
rect 7477 67408 7785 67428
rect 9588 67244 9640 67250
rect 9588 67186 9640 67192
rect 9109 66940 9417 66960
rect 9109 66938 9115 66940
rect 9171 66938 9195 66940
rect 9251 66938 9275 66940
rect 9331 66938 9355 66940
rect 9411 66938 9417 66940
rect 9171 66886 9173 66938
rect 9353 66886 9355 66938
rect 9109 66884 9115 66886
rect 9171 66884 9195 66886
rect 9251 66884 9275 66886
rect 9331 66884 9355 66886
rect 9411 66884 9417 66886
rect 9109 66864 9417 66884
rect 7477 66396 7785 66416
rect 7477 66394 7483 66396
rect 7539 66394 7563 66396
rect 7619 66394 7643 66396
rect 7699 66394 7723 66396
rect 7779 66394 7785 66396
rect 7539 66342 7541 66394
rect 7721 66342 7723 66394
rect 7477 66340 7483 66342
rect 7539 66340 7563 66342
rect 7619 66340 7643 66342
rect 7699 66340 7723 66342
rect 7779 66340 7785 66342
rect 7477 66320 7785 66340
rect 9109 65852 9417 65872
rect 9109 65850 9115 65852
rect 9171 65850 9195 65852
rect 9251 65850 9275 65852
rect 9331 65850 9355 65852
rect 9411 65850 9417 65852
rect 9171 65798 9173 65850
rect 9353 65798 9355 65850
rect 9109 65796 9115 65798
rect 9171 65796 9195 65798
rect 9251 65796 9275 65798
rect 9331 65796 9355 65798
rect 9411 65796 9417 65798
rect 9109 65776 9417 65796
rect 7477 65308 7785 65328
rect 7477 65306 7483 65308
rect 7539 65306 7563 65308
rect 7619 65306 7643 65308
rect 7699 65306 7723 65308
rect 7779 65306 7785 65308
rect 7539 65254 7541 65306
rect 7721 65254 7723 65306
rect 7477 65252 7483 65254
rect 7539 65252 7563 65254
rect 7619 65252 7643 65254
rect 7699 65252 7723 65254
rect 7779 65252 7785 65254
rect 7477 65232 7785 65252
rect 9600 65210 9628 67186
rect 9680 66156 9732 66162
rect 9680 66098 9732 66104
rect 9588 65204 9640 65210
rect 9588 65146 9640 65152
rect 9109 64764 9417 64784
rect 9109 64762 9115 64764
rect 9171 64762 9195 64764
rect 9251 64762 9275 64764
rect 9331 64762 9355 64764
rect 9411 64762 9417 64764
rect 9171 64710 9173 64762
rect 9353 64710 9355 64762
rect 9109 64708 9115 64710
rect 9171 64708 9195 64710
rect 9251 64708 9275 64710
rect 9331 64708 9355 64710
rect 9411 64708 9417 64710
rect 9109 64688 9417 64708
rect 7196 64388 7248 64394
rect 7196 64330 7248 64336
rect 7104 46368 7156 46374
rect 7104 46310 7156 46316
rect 7012 38480 7064 38486
rect 7012 38422 7064 38428
rect 6932 31726 7052 31754
rect 7024 28694 7052 31726
rect 7012 28688 7064 28694
rect 7012 28630 7064 28636
rect 7116 24682 7144 46310
rect 7208 30394 7236 64330
rect 7477 64220 7785 64240
rect 7477 64218 7483 64220
rect 7539 64218 7563 64220
rect 7619 64218 7643 64220
rect 7699 64218 7723 64220
rect 7779 64218 7785 64220
rect 7539 64166 7541 64218
rect 7721 64166 7723 64218
rect 7477 64164 7483 64166
rect 7539 64164 7563 64166
rect 7619 64164 7643 64166
rect 7699 64164 7723 64166
rect 7779 64164 7785 64166
rect 7477 64144 7785 64164
rect 9692 64122 9720 66098
rect 9784 66094 9812 67662
rect 9876 66842 9904 68274
rect 10046 68232 10102 68241
rect 10046 68167 10048 68176
rect 10100 68167 10102 68176
rect 10048 68138 10100 68144
rect 10048 67584 10100 67590
rect 10048 67526 10100 67532
rect 10060 67425 10088 67526
rect 10046 67416 10102 67425
rect 10046 67351 10102 67360
rect 10048 67040 10100 67046
rect 10048 66982 10100 66988
rect 9864 66836 9916 66842
rect 9864 66778 9916 66784
rect 10060 66745 10088 66982
rect 10046 66736 10102 66745
rect 10046 66671 10102 66680
rect 9772 66088 9824 66094
rect 9772 66030 9824 66036
rect 10048 65952 10100 65958
rect 10046 65920 10048 65929
rect 10100 65920 10102 65929
rect 10046 65855 10102 65864
rect 9864 65544 9916 65550
rect 9864 65486 9916 65492
rect 9876 64598 9904 65486
rect 10048 65408 10100 65414
rect 10048 65350 10100 65356
rect 10060 65249 10088 65350
rect 10046 65240 10102 65249
rect 10046 65175 10102 65184
rect 9864 64592 9916 64598
rect 9864 64534 9916 64540
rect 9772 64456 9824 64462
rect 9772 64398 9824 64404
rect 10046 64424 10102 64433
rect 9680 64116 9732 64122
rect 9680 64058 9732 64064
rect 8392 64048 8444 64054
rect 8392 63990 8444 63996
rect 8300 63776 8352 63782
rect 8300 63718 8352 63724
rect 7477 63132 7785 63152
rect 7477 63130 7483 63132
rect 7539 63130 7563 63132
rect 7619 63130 7643 63132
rect 7699 63130 7723 63132
rect 7779 63130 7785 63132
rect 7539 63078 7541 63130
rect 7721 63078 7723 63130
rect 7477 63076 7483 63078
rect 7539 63076 7563 63078
rect 7619 63076 7643 63078
rect 7699 63076 7723 63078
rect 7779 63076 7785 63078
rect 7477 63056 7785 63076
rect 7477 62044 7785 62064
rect 7477 62042 7483 62044
rect 7539 62042 7563 62044
rect 7619 62042 7643 62044
rect 7699 62042 7723 62044
rect 7779 62042 7785 62044
rect 7539 61990 7541 62042
rect 7721 61990 7723 62042
rect 7477 61988 7483 61990
rect 7539 61988 7563 61990
rect 7619 61988 7643 61990
rect 7699 61988 7723 61990
rect 7779 61988 7785 61990
rect 7477 61968 7785 61988
rect 7477 60956 7785 60976
rect 7477 60954 7483 60956
rect 7539 60954 7563 60956
rect 7619 60954 7643 60956
rect 7699 60954 7723 60956
rect 7779 60954 7785 60956
rect 7539 60902 7541 60954
rect 7721 60902 7723 60954
rect 7477 60900 7483 60902
rect 7539 60900 7563 60902
rect 7619 60900 7643 60902
rect 7699 60900 7723 60902
rect 7779 60900 7785 60902
rect 7477 60880 7785 60900
rect 7477 59868 7785 59888
rect 7477 59866 7483 59868
rect 7539 59866 7563 59868
rect 7619 59866 7643 59868
rect 7699 59866 7723 59868
rect 7779 59866 7785 59868
rect 7539 59814 7541 59866
rect 7721 59814 7723 59866
rect 7477 59812 7483 59814
rect 7539 59812 7563 59814
rect 7619 59812 7643 59814
rect 7699 59812 7723 59814
rect 7779 59812 7785 59814
rect 7477 59792 7785 59812
rect 7477 58780 7785 58800
rect 7477 58778 7483 58780
rect 7539 58778 7563 58780
rect 7619 58778 7643 58780
rect 7699 58778 7723 58780
rect 7779 58778 7785 58780
rect 7539 58726 7541 58778
rect 7721 58726 7723 58778
rect 7477 58724 7483 58726
rect 7539 58724 7563 58726
rect 7619 58724 7643 58726
rect 7699 58724 7723 58726
rect 7779 58724 7785 58726
rect 7477 58704 7785 58724
rect 7477 57692 7785 57712
rect 7477 57690 7483 57692
rect 7539 57690 7563 57692
rect 7619 57690 7643 57692
rect 7699 57690 7723 57692
rect 7779 57690 7785 57692
rect 7539 57638 7541 57690
rect 7721 57638 7723 57690
rect 7477 57636 7483 57638
rect 7539 57636 7563 57638
rect 7619 57636 7643 57638
rect 7699 57636 7723 57638
rect 7779 57636 7785 57638
rect 7477 57616 7785 57636
rect 7380 57384 7432 57390
rect 7380 57326 7432 57332
rect 7288 56908 7340 56914
rect 7288 56850 7340 56856
rect 7196 30388 7248 30394
rect 7196 30330 7248 30336
rect 7300 25498 7328 56850
rect 7392 46374 7420 57326
rect 7477 56604 7785 56624
rect 7477 56602 7483 56604
rect 7539 56602 7563 56604
rect 7619 56602 7643 56604
rect 7699 56602 7723 56604
rect 7779 56602 7785 56604
rect 7539 56550 7541 56602
rect 7721 56550 7723 56602
rect 7477 56548 7483 56550
rect 7539 56548 7563 56550
rect 7619 56548 7643 56550
rect 7699 56548 7723 56550
rect 7779 56548 7785 56550
rect 7477 56528 7785 56548
rect 7477 55516 7785 55536
rect 7477 55514 7483 55516
rect 7539 55514 7563 55516
rect 7619 55514 7643 55516
rect 7699 55514 7723 55516
rect 7779 55514 7785 55516
rect 7539 55462 7541 55514
rect 7721 55462 7723 55514
rect 7477 55460 7483 55462
rect 7539 55460 7563 55462
rect 7619 55460 7643 55462
rect 7699 55460 7723 55462
rect 7779 55460 7785 55462
rect 7477 55440 7785 55460
rect 7477 54428 7785 54448
rect 7477 54426 7483 54428
rect 7539 54426 7563 54428
rect 7619 54426 7643 54428
rect 7699 54426 7723 54428
rect 7779 54426 7785 54428
rect 7539 54374 7541 54426
rect 7721 54374 7723 54426
rect 7477 54372 7483 54374
rect 7539 54372 7563 54374
rect 7619 54372 7643 54374
rect 7699 54372 7723 54374
rect 7779 54372 7785 54374
rect 7477 54352 7785 54372
rect 7477 53340 7785 53360
rect 7477 53338 7483 53340
rect 7539 53338 7563 53340
rect 7619 53338 7643 53340
rect 7699 53338 7723 53340
rect 7779 53338 7785 53340
rect 7539 53286 7541 53338
rect 7721 53286 7723 53338
rect 7477 53284 7483 53286
rect 7539 53284 7563 53286
rect 7619 53284 7643 53286
rect 7699 53284 7723 53286
rect 7779 53284 7785 53286
rect 7477 53264 7785 53284
rect 7477 52252 7785 52272
rect 7477 52250 7483 52252
rect 7539 52250 7563 52252
rect 7619 52250 7643 52252
rect 7699 52250 7723 52252
rect 7779 52250 7785 52252
rect 7539 52198 7541 52250
rect 7721 52198 7723 52250
rect 7477 52196 7483 52198
rect 7539 52196 7563 52198
rect 7619 52196 7643 52198
rect 7699 52196 7723 52198
rect 7779 52196 7785 52198
rect 7477 52176 7785 52196
rect 8024 52080 8076 52086
rect 8024 52022 8076 52028
rect 7838 51504 7894 51513
rect 7838 51439 7894 51448
rect 7477 51164 7785 51184
rect 7477 51162 7483 51164
rect 7539 51162 7563 51164
rect 7619 51162 7643 51164
rect 7699 51162 7723 51164
rect 7779 51162 7785 51164
rect 7539 51110 7541 51162
rect 7721 51110 7723 51162
rect 7477 51108 7483 51110
rect 7539 51108 7563 51110
rect 7619 51108 7643 51110
rect 7699 51108 7723 51110
rect 7779 51108 7785 51110
rect 7477 51088 7785 51108
rect 7477 50076 7785 50096
rect 7477 50074 7483 50076
rect 7539 50074 7563 50076
rect 7619 50074 7643 50076
rect 7699 50074 7723 50076
rect 7779 50074 7785 50076
rect 7539 50022 7541 50074
rect 7721 50022 7723 50074
rect 7477 50020 7483 50022
rect 7539 50020 7563 50022
rect 7619 50020 7643 50022
rect 7699 50020 7723 50022
rect 7779 50020 7785 50022
rect 7477 50000 7785 50020
rect 7477 48988 7785 49008
rect 7477 48986 7483 48988
rect 7539 48986 7563 48988
rect 7619 48986 7643 48988
rect 7699 48986 7723 48988
rect 7779 48986 7785 48988
rect 7539 48934 7541 48986
rect 7721 48934 7723 48986
rect 7477 48932 7483 48934
rect 7539 48932 7563 48934
rect 7619 48932 7643 48934
rect 7699 48932 7723 48934
rect 7779 48932 7785 48934
rect 7477 48912 7785 48932
rect 7477 47900 7785 47920
rect 7477 47898 7483 47900
rect 7539 47898 7563 47900
rect 7619 47898 7643 47900
rect 7699 47898 7723 47900
rect 7779 47898 7785 47900
rect 7539 47846 7541 47898
rect 7721 47846 7723 47898
rect 7477 47844 7483 47846
rect 7539 47844 7563 47846
rect 7619 47844 7643 47846
rect 7699 47844 7723 47846
rect 7779 47844 7785 47846
rect 7477 47824 7785 47844
rect 7477 46812 7785 46832
rect 7477 46810 7483 46812
rect 7539 46810 7563 46812
rect 7619 46810 7643 46812
rect 7699 46810 7723 46812
rect 7779 46810 7785 46812
rect 7539 46758 7541 46810
rect 7721 46758 7723 46810
rect 7477 46756 7483 46758
rect 7539 46756 7563 46758
rect 7619 46756 7643 46758
rect 7699 46756 7723 46758
rect 7779 46756 7785 46758
rect 7477 46736 7785 46756
rect 7380 46368 7432 46374
rect 7380 46310 7432 46316
rect 7852 46186 7880 51439
rect 7932 46436 7984 46442
rect 7932 46378 7984 46384
rect 7392 46158 7880 46186
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 7104 24676 7156 24682
rect 7104 24618 7156 24624
rect 7392 22778 7420 46158
rect 7840 46096 7892 46102
rect 7840 46038 7892 46044
rect 7477 45724 7785 45744
rect 7477 45722 7483 45724
rect 7539 45722 7563 45724
rect 7619 45722 7643 45724
rect 7699 45722 7723 45724
rect 7779 45722 7785 45724
rect 7539 45670 7541 45722
rect 7721 45670 7723 45722
rect 7477 45668 7483 45670
rect 7539 45668 7563 45670
rect 7619 45668 7643 45670
rect 7699 45668 7723 45670
rect 7779 45668 7785 45670
rect 7477 45648 7785 45668
rect 7477 44636 7785 44656
rect 7477 44634 7483 44636
rect 7539 44634 7563 44636
rect 7619 44634 7643 44636
rect 7699 44634 7723 44636
rect 7779 44634 7785 44636
rect 7539 44582 7541 44634
rect 7721 44582 7723 44634
rect 7477 44580 7483 44582
rect 7539 44580 7563 44582
rect 7619 44580 7643 44582
rect 7699 44580 7723 44582
rect 7779 44580 7785 44582
rect 7477 44560 7785 44580
rect 7477 43548 7785 43568
rect 7477 43546 7483 43548
rect 7539 43546 7563 43548
rect 7619 43546 7643 43548
rect 7699 43546 7723 43548
rect 7779 43546 7785 43548
rect 7539 43494 7541 43546
rect 7721 43494 7723 43546
rect 7477 43492 7483 43494
rect 7539 43492 7563 43494
rect 7619 43492 7643 43494
rect 7699 43492 7723 43494
rect 7779 43492 7785 43494
rect 7477 43472 7785 43492
rect 7477 42460 7785 42480
rect 7477 42458 7483 42460
rect 7539 42458 7563 42460
rect 7619 42458 7643 42460
rect 7699 42458 7723 42460
rect 7779 42458 7785 42460
rect 7539 42406 7541 42458
rect 7721 42406 7723 42458
rect 7477 42404 7483 42406
rect 7539 42404 7563 42406
rect 7619 42404 7643 42406
rect 7699 42404 7723 42406
rect 7779 42404 7785 42406
rect 7477 42384 7785 42404
rect 7477 41372 7785 41392
rect 7477 41370 7483 41372
rect 7539 41370 7563 41372
rect 7619 41370 7643 41372
rect 7699 41370 7723 41372
rect 7779 41370 7785 41372
rect 7539 41318 7541 41370
rect 7721 41318 7723 41370
rect 7477 41316 7483 41318
rect 7539 41316 7563 41318
rect 7619 41316 7643 41318
rect 7699 41316 7723 41318
rect 7779 41316 7785 41318
rect 7477 41296 7785 41316
rect 7477 40284 7785 40304
rect 7477 40282 7483 40284
rect 7539 40282 7563 40284
rect 7619 40282 7643 40284
rect 7699 40282 7723 40284
rect 7779 40282 7785 40284
rect 7539 40230 7541 40282
rect 7721 40230 7723 40282
rect 7477 40228 7483 40230
rect 7539 40228 7563 40230
rect 7619 40228 7643 40230
rect 7699 40228 7723 40230
rect 7779 40228 7785 40230
rect 7477 40208 7785 40228
rect 7477 39196 7785 39216
rect 7477 39194 7483 39196
rect 7539 39194 7563 39196
rect 7619 39194 7643 39196
rect 7699 39194 7723 39196
rect 7779 39194 7785 39196
rect 7539 39142 7541 39194
rect 7721 39142 7723 39194
rect 7477 39140 7483 39142
rect 7539 39140 7563 39142
rect 7619 39140 7643 39142
rect 7699 39140 7723 39142
rect 7779 39140 7785 39142
rect 7477 39120 7785 39140
rect 7477 38108 7785 38128
rect 7477 38106 7483 38108
rect 7539 38106 7563 38108
rect 7619 38106 7643 38108
rect 7699 38106 7723 38108
rect 7779 38106 7785 38108
rect 7539 38054 7541 38106
rect 7721 38054 7723 38106
rect 7477 38052 7483 38054
rect 7539 38052 7563 38054
rect 7619 38052 7643 38054
rect 7699 38052 7723 38054
rect 7779 38052 7785 38054
rect 7477 38032 7785 38052
rect 7477 37020 7785 37040
rect 7477 37018 7483 37020
rect 7539 37018 7563 37020
rect 7619 37018 7643 37020
rect 7699 37018 7723 37020
rect 7779 37018 7785 37020
rect 7539 36966 7541 37018
rect 7721 36966 7723 37018
rect 7477 36964 7483 36966
rect 7539 36964 7563 36966
rect 7619 36964 7643 36966
rect 7699 36964 7723 36966
rect 7779 36964 7785 36966
rect 7477 36944 7785 36964
rect 7477 35932 7785 35952
rect 7477 35930 7483 35932
rect 7539 35930 7563 35932
rect 7619 35930 7643 35932
rect 7699 35930 7723 35932
rect 7779 35930 7785 35932
rect 7539 35878 7541 35930
rect 7721 35878 7723 35930
rect 7477 35876 7483 35878
rect 7539 35876 7563 35878
rect 7619 35876 7643 35878
rect 7699 35876 7723 35878
rect 7779 35876 7785 35878
rect 7477 35856 7785 35876
rect 7477 34844 7785 34864
rect 7477 34842 7483 34844
rect 7539 34842 7563 34844
rect 7619 34842 7643 34844
rect 7699 34842 7723 34844
rect 7779 34842 7785 34844
rect 7539 34790 7541 34842
rect 7721 34790 7723 34842
rect 7477 34788 7483 34790
rect 7539 34788 7563 34790
rect 7619 34788 7643 34790
rect 7699 34788 7723 34790
rect 7779 34788 7785 34790
rect 7477 34768 7785 34788
rect 7477 33756 7785 33776
rect 7477 33754 7483 33756
rect 7539 33754 7563 33756
rect 7619 33754 7643 33756
rect 7699 33754 7723 33756
rect 7779 33754 7785 33756
rect 7539 33702 7541 33754
rect 7721 33702 7723 33754
rect 7477 33700 7483 33702
rect 7539 33700 7563 33702
rect 7619 33700 7643 33702
rect 7699 33700 7723 33702
rect 7779 33700 7785 33702
rect 7477 33680 7785 33700
rect 7477 32668 7785 32688
rect 7477 32666 7483 32668
rect 7539 32666 7563 32668
rect 7619 32666 7643 32668
rect 7699 32666 7723 32668
rect 7779 32666 7785 32668
rect 7539 32614 7541 32666
rect 7721 32614 7723 32666
rect 7477 32612 7483 32614
rect 7539 32612 7563 32614
rect 7619 32612 7643 32614
rect 7699 32612 7723 32614
rect 7779 32612 7785 32614
rect 7477 32592 7785 32612
rect 7477 31580 7785 31600
rect 7477 31578 7483 31580
rect 7539 31578 7563 31580
rect 7619 31578 7643 31580
rect 7699 31578 7723 31580
rect 7779 31578 7785 31580
rect 7539 31526 7541 31578
rect 7721 31526 7723 31578
rect 7477 31524 7483 31526
rect 7539 31524 7563 31526
rect 7619 31524 7643 31526
rect 7699 31524 7723 31526
rect 7779 31524 7785 31526
rect 7477 31504 7785 31524
rect 7477 30492 7785 30512
rect 7477 30490 7483 30492
rect 7539 30490 7563 30492
rect 7619 30490 7643 30492
rect 7699 30490 7723 30492
rect 7779 30490 7785 30492
rect 7539 30438 7541 30490
rect 7721 30438 7723 30490
rect 7477 30436 7483 30438
rect 7539 30436 7563 30438
rect 7619 30436 7643 30438
rect 7699 30436 7723 30438
rect 7779 30436 7785 30438
rect 7477 30416 7785 30436
rect 7477 29404 7785 29424
rect 7477 29402 7483 29404
rect 7539 29402 7563 29404
rect 7619 29402 7643 29404
rect 7699 29402 7723 29404
rect 7779 29402 7785 29404
rect 7539 29350 7541 29402
rect 7721 29350 7723 29402
rect 7477 29348 7483 29350
rect 7539 29348 7563 29350
rect 7619 29348 7643 29350
rect 7699 29348 7723 29350
rect 7779 29348 7785 29350
rect 7477 29328 7785 29348
rect 7477 28316 7785 28336
rect 7477 28314 7483 28316
rect 7539 28314 7563 28316
rect 7619 28314 7643 28316
rect 7699 28314 7723 28316
rect 7779 28314 7785 28316
rect 7539 28262 7541 28314
rect 7721 28262 7723 28314
rect 7477 28260 7483 28262
rect 7539 28260 7563 28262
rect 7619 28260 7643 28262
rect 7699 28260 7723 28262
rect 7779 28260 7785 28262
rect 7477 28240 7785 28260
rect 7477 27228 7785 27248
rect 7477 27226 7483 27228
rect 7539 27226 7563 27228
rect 7619 27226 7643 27228
rect 7699 27226 7723 27228
rect 7779 27226 7785 27228
rect 7539 27174 7541 27226
rect 7721 27174 7723 27226
rect 7477 27172 7483 27174
rect 7539 27172 7563 27174
rect 7619 27172 7643 27174
rect 7699 27172 7723 27174
rect 7779 27172 7785 27174
rect 7477 27152 7785 27172
rect 7477 26140 7785 26160
rect 7477 26138 7483 26140
rect 7539 26138 7563 26140
rect 7619 26138 7643 26140
rect 7699 26138 7723 26140
rect 7779 26138 7785 26140
rect 7539 26086 7541 26138
rect 7721 26086 7723 26138
rect 7477 26084 7483 26086
rect 7539 26084 7563 26086
rect 7619 26084 7643 26086
rect 7699 26084 7723 26086
rect 7779 26084 7785 26086
rect 7477 26064 7785 26084
rect 7477 25052 7785 25072
rect 7477 25050 7483 25052
rect 7539 25050 7563 25052
rect 7619 25050 7643 25052
rect 7699 25050 7723 25052
rect 7779 25050 7785 25052
rect 7539 24998 7541 25050
rect 7721 24998 7723 25050
rect 7477 24996 7483 24998
rect 7539 24996 7563 24998
rect 7619 24996 7643 24998
rect 7699 24996 7723 24998
rect 7779 24996 7785 24998
rect 7477 24976 7785 24996
rect 7477 23964 7785 23984
rect 7477 23962 7483 23964
rect 7539 23962 7563 23964
rect 7619 23962 7643 23964
rect 7699 23962 7723 23964
rect 7779 23962 7785 23964
rect 7539 23910 7541 23962
rect 7721 23910 7723 23962
rect 7477 23908 7483 23910
rect 7539 23908 7563 23910
rect 7619 23908 7643 23910
rect 7699 23908 7723 23910
rect 7779 23908 7785 23910
rect 7477 23888 7785 23908
rect 7852 23322 7880 46038
rect 7840 23316 7892 23322
rect 7840 23258 7892 23264
rect 7477 22876 7785 22896
rect 7477 22874 7483 22876
rect 7539 22874 7563 22876
rect 7619 22874 7643 22876
rect 7699 22874 7723 22876
rect 7779 22874 7785 22876
rect 7539 22822 7541 22874
rect 7721 22822 7723 22874
rect 7477 22820 7483 22822
rect 7539 22820 7563 22822
rect 7619 22820 7643 22822
rect 7699 22820 7723 22822
rect 7779 22820 7785 22822
rect 7477 22800 7785 22820
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7477 21788 7785 21808
rect 7477 21786 7483 21788
rect 7539 21786 7563 21788
rect 7619 21786 7643 21788
rect 7699 21786 7723 21788
rect 7779 21786 7785 21788
rect 7539 21734 7541 21786
rect 7721 21734 7723 21786
rect 7477 21732 7483 21734
rect 7539 21732 7563 21734
rect 7619 21732 7643 21734
rect 7699 21732 7723 21734
rect 7779 21732 7785 21734
rect 7477 21712 7785 21732
rect 7477 20700 7785 20720
rect 7477 20698 7483 20700
rect 7539 20698 7563 20700
rect 7619 20698 7643 20700
rect 7699 20698 7723 20700
rect 7779 20698 7785 20700
rect 7539 20646 7541 20698
rect 7721 20646 7723 20698
rect 7477 20644 7483 20646
rect 7539 20644 7563 20646
rect 7619 20644 7643 20646
rect 7699 20644 7723 20646
rect 7779 20644 7785 20646
rect 7477 20624 7785 20644
rect 7477 19612 7785 19632
rect 7477 19610 7483 19612
rect 7539 19610 7563 19612
rect 7619 19610 7643 19612
rect 7699 19610 7723 19612
rect 7779 19610 7785 19612
rect 7539 19558 7541 19610
rect 7721 19558 7723 19610
rect 7477 19556 7483 19558
rect 7539 19556 7563 19558
rect 7619 19556 7643 19558
rect 7699 19556 7723 19558
rect 7779 19556 7785 19558
rect 7477 19536 7785 19556
rect 7477 18524 7785 18544
rect 7477 18522 7483 18524
rect 7539 18522 7563 18524
rect 7619 18522 7643 18524
rect 7699 18522 7723 18524
rect 7779 18522 7785 18524
rect 7539 18470 7541 18522
rect 7721 18470 7723 18522
rect 7477 18468 7483 18470
rect 7539 18468 7563 18470
rect 7619 18468 7643 18470
rect 7699 18468 7723 18470
rect 7779 18468 7785 18470
rect 7477 18448 7785 18468
rect 7944 17678 7972 46378
rect 8036 22098 8064 52022
rect 8116 50516 8168 50522
rect 8116 50458 8168 50464
rect 8128 46102 8156 50458
rect 8116 46096 8168 46102
rect 8116 46038 8168 46044
rect 8312 29510 8340 63718
rect 8404 31210 8432 63990
rect 9784 63850 9812 64398
rect 10046 64359 10102 64368
rect 10060 64326 10088 64359
rect 10048 64320 10100 64326
rect 10048 64262 10100 64268
rect 9864 63980 9916 63986
rect 9864 63922 9916 63928
rect 9772 63844 9824 63850
rect 9772 63786 9824 63792
rect 9109 63676 9417 63696
rect 9109 63674 9115 63676
rect 9171 63674 9195 63676
rect 9251 63674 9275 63676
rect 9331 63674 9355 63676
rect 9411 63674 9417 63676
rect 9171 63622 9173 63674
rect 9353 63622 9355 63674
rect 9109 63620 9115 63622
rect 9171 63620 9195 63622
rect 9251 63620 9275 63622
rect 9331 63620 9355 63622
rect 9411 63620 9417 63622
rect 9109 63600 9417 63620
rect 9876 63510 9904 63922
rect 10048 63776 10100 63782
rect 10048 63718 10100 63724
rect 10060 63617 10088 63718
rect 10046 63608 10102 63617
rect 10046 63543 10102 63552
rect 9864 63504 9916 63510
rect 9864 63446 9916 63452
rect 9864 63368 9916 63374
rect 9864 63310 9916 63316
rect 8484 62756 8536 62762
rect 8484 62698 8536 62704
rect 8392 31204 8444 31210
rect 8392 31146 8444 31152
rect 8496 29850 8524 62698
rect 9876 62694 9904 63310
rect 10048 63232 10100 63238
rect 10048 63174 10100 63180
rect 10060 62937 10088 63174
rect 10046 62928 10102 62937
rect 10046 62863 10102 62872
rect 9864 62688 9916 62694
rect 9864 62630 9916 62636
rect 9109 62588 9417 62608
rect 9109 62586 9115 62588
rect 9171 62586 9195 62588
rect 9251 62586 9275 62588
rect 9331 62586 9355 62588
rect 9411 62586 9417 62588
rect 9171 62534 9173 62586
rect 9353 62534 9355 62586
rect 9109 62532 9115 62534
rect 9171 62532 9195 62534
rect 9251 62532 9275 62534
rect 9331 62532 9355 62534
rect 9411 62532 9417 62534
rect 9109 62512 9417 62532
rect 10048 62144 10100 62150
rect 10046 62112 10048 62121
rect 10100 62112 10102 62121
rect 10046 62047 10102 62056
rect 10048 61600 10100 61606
rect 10048 61542 10100 61548
rect 9109 61500 9417 61520
rect 9109 61498 9115 61500
rect 9171 61498 9195 61500
rect 9251 61498 9275 61500
rect 9331 61498 9355 61500
rect 9411 61498 9417 61500
rect 9171 61446 9173 61498
rect 9353 61446 9355 61498
rect 9109 61444 9115 61446
rect 9171 61444 9195 61446
rect 9251 61444 9275 61446
rect 9331 61444 9355 61446
rect 9411 61444 9417 61446
rect 9109 61424 9417 61444
rect 10060 61441 10088 61542
rect 10046 61432 10102 61441
rect 10046 61367 10102 61376
rect 10046 60616 10102 60625
rect 10046 60551 10048 60560
rect 10100 60551 10102 60560
rect 10048 60522 10100 60528
rect 9109 60412 9417 60432
rect 9109 60410 9115 60412
rect 9171 60410 9195 60412
rect 9251 60410 9275 60412
rect 9331 60410 9355 60412
rect 9411 60410 9417 60412
rect 9171 60358 9173 60410
rect 9353 60358 9355 60410
rect 9109 60356 9115 60358
rect 9171 60356 9195 60358
rect 9251 60356 9275 60358
rect 9331 60356 9355 60358
rect 9411 60356 9417 60358
rect 9109 60336 9417 60356
rect 9772 60104 9824 60110
rect 9772 60046 9824 60052
rect 9109 59324 9417 59344
rect 9109 59322 9115 59324
rect 9171 59322 9195 59324
rect 9251 59322 9275 59324
rect 9331 59322 9355 59324
rect 9411 59322 9417 59324
rect 9171 59270 9173 59322
rect 9353 59270 9355 59322
rect 9109 59268 9115 59270
rect 9171 59268 9195 59270
rect 9251 59268 9275 59270
rect 9331 59268 9355 59270
rect 9411 59268 9417 59270
rect 9109 59248 9417 59268
rect 9109 58236 9417 58256
rect 9109 58234 9115 58236
rect 9171 58234 9195 58236
rect 9251 58234 9275 58236
rect 9331 58234 9355 58236
rect 9411 58234 9417 58236
rect 9171 58182 9173 58234
rect 9353 58182 9355 58234
rect 9109 58180 9115 58182
rect 9171 58180 9195 58182
rect 9251 58180 9275 58182
rect 9331 58180 9355 58182
rect 9411 58180 9417 58182
rect 9109 58160 9417 58180
rect 8576 57860 8628 57866
rect 8576 57802 8628 57808
rect 8484 29844 8536 29850
rect 8484 29786 8536 29792
rect 8300 29504 8352 29510
rect 8300 29446 8352 29452
rect 8588 26042 8616 57802
rect 9109 57148 9417 57168
rect 9109 57146 9115 57148
rect 9171 57146 9195 57148
rect 9251 57146 9275 57148
rect 9331 57146 9355 57148
rect 9411 57146 9417 57148
rect 9171 57094 9173 57146
rect 9353 57094 9355 57146
rect 9109 57092 9115 57094
rect 9171 57092 9195 57094
rect 9251 57092 9275 57094
rect 9331 57092 9355 57094
rect 9411 57092 9417 57094
rect 9109 57072 9417 57092
rect 9784 56982 9812 60046
rect 10048 59968 10100 59974
rect 10046 59936 10048 59945
rect 10100 59936 10102 59945
rect 10046 59871 10102 59880
rect 9864 59628 9916 59634
rect 9864 59570 9916 59576
rect 9876 57322 9904 59570
rect 10048 59424 10100 59430
rect 10048 59366 10100 59372
rect 10060 59129 10088 59366
rect 10046 59120 10102 59129
rect 10046 59055 10102 59064
rect 10046 58440 10102 58449
rect 10046 58375 10048 58384
rect 10100 58375 10102 58384
rect 10048 58346 10100 58352
rect 10048 57792 10100 57798
rect 10048 57734 10100 57740
rect 10060 57633 10088 57734
rect 10046 57624 10102 57633
rect 10046 57559 10102 57568
rect 9864 57316 9916 57322
rect 9864 57258 9916 57264
rect 10048 57248 10100 57254
rect 10048 57190 10100 57196
rect 9772 56976 9824 56982
rect 10060 56953 10088 57190
rect 9772 56918 9824 56924
rect 10046 56944 10102 56953
rect 10046 56879 10102 56888
rect 8668 56228 8720 56234
rect 8668 56170 8720 56176
rect 8680 26586 8708 56170
rect 10048 56160 10100 56166
rect 10046 56128 10048 56137
rect 10100 56128 10102 56137
rect 9109 56060 9417 56080
rect 10046 56063 10102 56072
rect 9109 56058 9115 56060
rect 9171 56058 9195 56060
rect 9251 56058 9275 56060
rect 9331 56058 9355 56060
rect 9411 56058 9417 56060
rect 9171 56006 9173 56058
rect 9353 56006 9355 56058
rect 9109 56004 9115 56006
rect 9171 56004 9195 56006
rect 9251 56004 9275 56006
rect 9331 56004 9355 56006
rect 9411 56004 9417 56006
rect 9109 55984 9417 56004
rect 10048 55616 10100 55622
rect 10048 55558 10100 55564
rect 10060 55321 10088 55558
rect 10046 55312 10102 55321
rect 8760 55276 8812 55282
rect 10046 55247 10102 55256
rect 8760 55218 8812 55224
rect 8772 28422 8800 55218
rect 9109 54972 9417 54992
rect 9109 54970 9115 54972
rect 9171 54970 9195 54972
rect 9251 54970 9275 54972
rect 9331 54970 9355 54972
rect 9411 54970 9417 54972
rect 9171 54918 9173 54970
rect 9353 54918 9355 54970
rect 9109 54916 9115 54918
rect 9171 54916 9195 54918
rect 9251 54916 9275 54918
rect 9331 54916 9355 54918
rect 9411 54916 9417 54918
rect 9109 54896 9417 54916
rect 10140 54664 10192 54670
rect 10138 54632 10140 54641
rect 10192 54632 10194 54641
rect 10138 54567 10194 54576
rect 9956 54528 10008 54534
rect 9956 54470 10008 54476
rect 9864 53984 9916 53990
rect 9864 53926 9916 53932
rect 9109 53884 9417 53904
rect 9109 53882 9115 53884
rect 9171 53882 9195 53884
rect 9251 53882 9275 53884
rect 9331 53882 9355 53884
rect 9411 53882 9417 53884
rect 9171 53830 9173 53882
rect 9353 53830 9355 53882
rect 9109 53828 9115 53830
rect 9171 53828 9195 53830
rect 9251 53828 9275 53830
rect 9331 53828 9355 53830
rect 9411 53828 9417 53830
rect 9109 53808 9417 53828
rect 9876 53106 9904 53926
rect 9968 53582 9996 54470
rect 10140 54188 10192 54194
rect 10140 54130 10192 54136
rect 10152 53825 10180 54130
rect 10138 53816 10194 53825
rect 10138 53751 10194 53760
rect 9956 53576 10008 53582
rect 9956 53518 10008 53524
rect 10140 53576 10192 53582
rect 10140 53518 10192 53524
rect 9956 53440 10008 53446
rect 9956 53382 10008 53388
rect 9864 53100 9916 53106
rect 9864 53042 9916 53048
rect 9109 52796 9417 52816
rect 9109 52794 9115 52796
rect 9171 52794 9195 52796
rect 9251 52794 9275 52796
rect 9331 52794 9355 52796
rect 9411 52794 9417 52796
rect 9171 52742 9173 52794
rect 9353 52742 9355 52794
rect 9109 52740 9115 52742
rect 9171 52740 9195 52742
rect 9251 52740 9275 52742
rect 9331 52740 9355 52742
rect 9411 52740 9417 52742
rect 9109 52720 9417 52740
rect 9968 52494 9996 53382
rect 10152 53145 10180 53518
rect 10138 53136 10194 53145
rect 10138 53071 10194 53080
rect 9956 52488 10008 52494
rect 9956 52430 10008 52436
rect 10140 52488 10192 52494
rect 10140 52430 10192 52436
rect 9496 52352 9548 52358
rect 10152 52329 10180 52430
rect 9496 52294 9548 52300
rect 10138 52320 10194 52329
rect 9109 51708 9417 51728
rect 9109 51706 9115 51708
rect 9171 51706 9195 51708
rect 9251 51706 9275 51708
rect 9331 51706 9355 51708
rect 9411 51706 9417 51708
rect 9171 51654 9173 51706
rect 9353 51654 9355 51706
rect 9109 51652 9115 51654
rect 9171 51652 9195 51654
rect 9251 51652 9275 51654
rect 9331 51652 9355 51654
rect 9411 51652 9417 51654
rect 9109 51632 9417 51652
rect 9508 51406 9536 52294
rect 10138 52255 10194 52264
rect 10140 52012 10192 52018
rect 10140 51954 10192 51960
rect 9956 51808 10008 51814
rect 9956 51750 10008 51756
rect 9496 51400 9548 51406
rect 9496 51342 9548 51348
rect 9968 51066 9996 51750
rect 10152 51649 10180 51954
rect 10138 51640 10194 51649
rect 10138 51575 10194 51584
rect 9956 51060 10008 51066
rect 9956 51002 10008 51008
rect 10140 50924 10192 50930
rect 10140 50866 10192 50872
rect 10152 50833 10180 50866
rect 10138 50824 10194 50833
rect 10138 50759 10194 50768
rect 9956 50720 10008 50726
rect 9956 50662 10008 50668
rect 9109 50620 9417 50640
rect 9109 50618 9115 50620
rect 9171 50618 9195 50620
rect 9251 50618 9275 50620
rect 9331 50618 9355 50620
rect 9411 50618 9417 50620
rect 9171 50566 9173 50618
rect 9353 50566 9355 50618
rect 9109 50564 9115 50566
rect 9171 50564 9195 50566
rect 9251 50564 9275 50566
rect 9331 50564 9355 50566
rect 9411 50564 9417 50566
rect 9109 50544 9417 50564
rect 9968 50318 9996 50662
rect 9956 50312 10008 50318
rect 9956 50254 10008 50260
rect 10140 50312 10192 50318
rect 10140 50254 10192 50260
rect 9956 50176 10008 50182
rect 10152 50153 10180 50254
rect 9956 50118 10008 50124
rect 10138 50144 10194 50153
rect 9968 49842 9996 50118
rect 10138 50079 10194 50088
rect 9956 49836 10008 49842
rect 9956 49778 10008 49784
rect 10140 49700 10192 49706
rect 10140 49642 10192 49648
rect 9109 49532 9417 49552
rect 9109 49530 9115 49532
rect 9171 49530 9195 49532
rect 9251 49530 9275 49532
rect 9331 49530 9355 49532
rect 9411 49530 9417 49532
rect 9171 49478 9173 49530
rect 9353 49478 9355 49530
rect 9109 49476 9115 49478
rect 9171 49476 9195 49478
rect 9251 49476 9275 49478
rect 9331 49476 9355 49478
rect 9411 49476 9417 49478
rect 9109 49456 9417 49476
rect 10152 49337 10180 49642
rect 10138 49328 10194 49337
rect 10138 49263 10194 49272
rect 10140 48748 10192 48754
rect 10140 48690 10192 48696
rect 10152 48657 10180 48690
rect 10138 48648 10194 48657
rect 10138 48583 10194 48592
rect 9956 48544 10008 48550
rect 9956 48486 10008 48492
rect 9109 48444 9417 48464
rect 9109 48442 9115 48444
rect 9171 48442 9195 48444
rect 9251 48442 9275 48444
rect 9331 48442 9355 48444
rect 9411 48442 9417 48444
rect 9171 48390 9173 48442
rect 9353 48390 9355 48442
rect 9109 48388 9115 48390
rect 9171 48388 9195 48390
rect 9251 48388 9275 48390
rect 9331 48388 9355 48390
rect 9411 48388 9417 48390
rect 9109 48368 9417 48388
rect 9864 48000 9916 48006
rect 9864 47942 9916 47948
rect 9109 47356 9417 47376
rect 9109 47354 9115 47356
rect 9171 47354 9195 47356
rect 9251 47354 9275 47356
rect 9331 47354 9355 47356
rect 9411 47354 9417 47356
rect 9171 47302 9173 47354
rect 9353 47302 9355 47354
rect 9109 47300 9115 47302
rect 9171 47300 9195 47302
rect 9251 47300 9275 47302
rect 9331 47300 9355 47302
rect 9411 47300 9417 47302
rect 9109 47280 9417 47300
rect 9876 46578 9904 47942
rect 9968 47666 9996 48486
rect 10140 48136 10192 48142
rect 10140 48078 10192 48084
rect 10152 47841 10180 48078
rect 10138 47832 10194 47841
rect 10138 47767 10194 47776
rect 9956 47660 10008 47666
rect 9956 47602 10008 47608
rect 10140 47048 10192 47054
rect 10138 47016 10140 47025
rect 10192 47016 10194 47025
rect 10138 46951 10194 46960
rect 9864 46572 9916 46578
rect 9864 46514 9916 46520
rect 10140 46572 10192 46578
rect 10140 46514 10192 46520
rect 9956 46368 10008 46374
rect 10152 46345 10180 46514
rect 9956 46310 10008 46316
rect 10138 46336 10194 46345
rect 9109 46268 9417 46288
rect 9109 46266 9115 46268
rect 9171 46266 9195 46268
rect 9251 46266 9275 46268
rect 9331 46266 9355 46268
rect 9411 46266 9417 46268
rect 9171 46214 9173 46266
rect 9353 46214 9355 46266
rect 9109 46212 9115 46214
rect 9171 46212 9195 46214
rect 9251 46212 9275 46214
rect 9331 46212 9355 46214
rect 9411 46212 9417 46214
rect 9109 46192 9417 46212
rect 9864 45824 9916 45830
rect 9864 45766 9916 45772
rect 9109 45180 9417 45200
rect 9109 45178 9115 45180
rect 9171 45178 9195 45180
rect 9251 45178 9275 45180
rect 9331 45178 9355 45180
rect 9411 45178 9417 45180
rect 9171 45126 9173 45178
rect 9353 45126 9355 45178
rect 9109 45124 9115 45126
rect 9171 45124 9195 45126
rect 9251 45124 9275 45126
rect 9331 45124 9355 45126
rect 9411 45124 9417 45126
rect 9109 45104 9417 45124
rect 9876 44878 9904 45766
rect 9968 45490 9996 46310
rect 10138 46271 10194 46280
rect 10140 45960 10192 45966
rect 10140 45902 10192 45908
rect 10152 45529 10180 45902
rect 10138 45520 10194 45529
rect 9956 45484 10008 45490
rect 10138 45455 10194 45464
rect 9956 45426 10008 45432
rect 9864 44872 9916 44878
rect 10140 44872 10192 44878
rect 9864 44814 9916 44820
rect 10138 44840 10140 44849
rect 10192 44840 10194 44849
rect 10138 44775 10194 44784
rect 9956 44736 10008 44742
rect 9956 44678 10008 44684
rect 9864 44192 9916 44198
rect 9864 44134 9916 44140
rect 9109 44092 9417 44112
rect 9109 44090 9115 44092
rect 9171 44090 9195 44092
rect 9251 44090 9275 44092
rect 9331 44090 9355 44092
rect 9411 44090 9417 44092
rect 9171 44038 9173 44090
rect 9353 44038 9355 44090
rect 9109 44036 9115 44038
rect 9171 44036 9195 44038
rect 9251 44036 9275 44038
rect 9331 44036 9355 44038
rect 9411 44036 9417 44038
rect 9109 44016 9417 44036
rect 9772 43648 9824 43654
rect 9772 43590 9824 43596
rect 9109 43004 9417 43024
rect 9109 43002 9115 43004
rect 9171 43002 9195 43004
rect 9251 43002 9275 43004
rect 9331 43002 9355 43004
rect 9411 43002 9417 43004
rect 9171 42950 9173 43002
rect 9353 42950 9355 43002
rect 9109 42948 9115 42950
rect 9171 42948 9195 42950
rect 9251 42948 9275 42950
rect 9331 42948 9355 42950
rect 9411 42948 9417 42950
rect 9109 42928 9417 42948
rect 9496 42696 9548 42702
rect 9496 42638 9548 42644
rect 9109 41916 9417 41936
rect 9109 41914 9115 41916
rect 9171 41914 9195 41916
rect 9251 41914 9275 41916
rect 9331 41914 9355 41916
rect 9411 41914 9417 41916
rect 9171 41862 9173 41914
rect 9353 41862 9355 41914
rect 9109 41860 9115 41862
rect 9171 41860 9195 41862
rect 9251 41860 9275 41862
rect 9331 41860 9355 41862
rect 9411 41860 9417 41862
rect 9109 41840 9417 41860
rect 9109 40828 9417 40848
rect 9109 40826 9115 40828
rect 9171 40826 9195 40828
rect 9251 40826 9275 40828
rect 9331 40826 9355 40828
rect 9411 40826 9417 40828
rect 9171 40774 9173 40826
rect 9353 40774 9355 40826
rect 9109 40772 9115 40774
rect 9171 40772 9195 40774
rect 9251 40772 9275 40774
rect 9331 40772 9355 40774
rect 9411 40772 9417 40774
rect 9109 40752 9417 40772
rect 9109 39740 9417 39760
rect 9109 39738 9115 39740
rect 9171 39738 9195 39740
rect 9251 39738 9275 39740
rect 9331 39738 9355 39740
rect 9411 39738 9417 39740
rect 9171 39686 9173 39738
rect 9353 39686 9355 39738
rect 9109 39684 9115 39686
rect 9171 39684 9195 39686
rect 9251 39684 9275 39686
rect 9331 39684 9355 39686
rect 9411 39684 9417 39686
rect 9109 39664 9417 39684
rect 9109 38652 9417 38672
rect 9109 38650 9115 38652
rect 9171 38650 9195 38652
rect 9251 38650 9275 38652
rect 9331 38650 9355 38652
rect 9411 38650 9417 38652
rect 9171 38598 9173 38650
rect 9353 38598 9355 38650
rect 9109 38596 9115 38598
rect 9171 38596 9195 38598
rect 9251 38596 9275 38598
rect 9331 38596 9355 38598
rect 9411 38596 9417 38598
rect 9109 38576 9417 38596
rect 9109 37564 9417 37584
rect 9109 37562 9115 37564
rect 9171 37562 9195 37564
rect 9251 37562 9275 37564
rect 9331 37562 9355 37564
rect 9411 37562 9417 37564
rect 9171 37510 9173 37562
rect 9353 37510 9355 37562
rect 9109 37508 9115 37510
rect 9171 37508 9195 37510
rect 9251 37508 9275 37510
rect 9331 37508 9355 37510
rect 9411 37508 9417 37510
rect 9109 37488 9417 37508
rect 9109 36476 9417 36496
rect 9109 36474 9115 36476
rect 9171 36474 9195 36476
rect 9251 36474 9275 36476
rect 9331 36474 9355 36476
rect 9411 36474 9417 36476
rect 9171 36422 9173 36474
rect 9353 36422 9355 36474
rect 9109 36420 9115 36422
rect 9171 36420 9195 36422
rect 9251 36420 9275 36422
rect 9331 36420 9355 36422
rect 9411 36420 9417 36422
rect 9109 36400 9417 36420
rect 9109 35388 9417 35408
rect 9109 35386 9115 35388
rect 9171 35386 9195 35388
rect 9251 35386 9275 35388
rect 9331 35386 9355 35388
rect 9411 35386 9417 35388
rect 9171 35334 9173 35386
rect 9353 35334 9355 35386
rect 9109 35332 9115 35334
rect 9171 35332 9195 35334
rect 9251 35332 9275 35334
rect 9331 35332 9355 35334
rect 9411 35332 9417 35334
rect 9109 35312 9417 35332
rect 9109 34300 9417 34320
rect 9109 34298 9115 34300
rect 9171 34298 9195 34300
rect 9251 34298 9275 34300
rect 9331 34298 9355 34300
rect 9411 34298 9417 34300
rect 9171 34246 9173 34298
rect 9353 34246 9355 34298
rect 9109 34244 9115 34246
rect 9171 34244 9195 34246
rect 9251 34244 9275 34246
rect 9331 34244 9355 34246
rect 9411 34244 9417 34246
rect 9109 34224 9417 34244
rect 9109 33212 9417 33232
rect 9109 33210 9115 33212
rect 9171 33210 9195 33212
rect 9251 33210 9275 33212
rect 9331 33210 9355 33212
rect 9411 33210 9417 33212
rect 9171 33158 9173 33210
rect 9353 33158 9355 33210
rect 9109 33156 9115 33158
rect 9171 33156 9195 33158
rect 9251 33156 9275 33158
rect 9331 33156 9355 33158
rect 9411 33156 9417 33158
rect 9109 33136 9417 33156
rect 9109 32124 9417 32144
rect 9109 32122 9115 32124
rect 9171 32122 9195 32124
rect 9251 32122 9275 32124
rect 9331 32122 9355 32124
rect 9411 32122 9417 32124
rect 9171 32070 9173 32122
rect 9353 32070 9355 32122
rect 9109 32068 9115 32070
rect 9171 32068 9195 32070
rect 9251 32068 9275 32070
rect 9331 32068 9355 32070
rect 9411 32068 9417 32070
rect 9109 32048 9417 32068
rect 9109 31036 9417 31056
rect 9109 31034 9115 31036
rect 9171 31034 9195 31036
rect 9251 31034 9275 31036
rect 9331 31034 9355 31036
rect 9411 31034 9417 31036
rect 9171 30982 9173 31034
rect 9353 30982 9355 31034
rect 9109 30980 9115 30982
rect 9171 30980 9195 30982
rect 9251 30980 9275 30982
rect 9331 30980 9355 30982
rect 9411 30980 9417 30982
rect 9109 30960 9417 30980
rect 9109 29948 9417 29968
rect 9109 29946 9115 29948
rect 9171 29946 9195 29948
rect 9251 29946 9275 29948
rect 9331 29946 9355 29948
rect 9411 29946 9417 29948
rect 9171 29894 9173 29946
rect 9353 29894 9355 29946
rect 9109 29892 9115 29894
rect 9171 29892 9195 29894
rect 9251 29892 9275 29894
rect 9331 29892 9355 29894
rect 9411 29892 9417 29894
rect 9109 29872 9417 29892
rect 9109 28860 9417 28880
rect 9109 28858 9115 28860
rect 9171 28858 9195 28860
rect 9251 28858 9275 28860
rect 9331 28858 9355 28860
rect 9411 28858 9417 28860
rect 9171 28806 9173 28858
rect 9353 28806 9355 28858
rect 9109 28804 9115 28806
rect 9171 28804 9195 28806
rect 9251 28804 9275 28806
rect 9331 28804 9355 28806
rect 9411 28804 9417 28806
rect 9109 28784 9417 28804
rect 8760 28416 8812 28422
rect 8760 28358 8812 28364
rect 9109 27772 9417 27792
rect 9109 27770 9115 27772
rect 9171 27770 9195 27772
rect 9251 27770 9275 27772
rect 9331 27770 9355 27772
rect 9411 27770 9417 27772
rect 9171 27718 9173 27770
rect 9353 27718 9355 27770
rect 9109 27716 9115 27718
rect 9171 27716 9195 27718
rect 9251 27716 9275 27718
rect 9331 27716 9355 27718
rect 9411 27716 9417 27718
rect 9109 27696 9417 27716
rect 9109 26684 9417 26704
rect 9109 26682 9115 26684
rect 9171 26682 9195 26684
rect 9251 26682 9275 26684
rect 9331 26682 9355 26684
rect 9411 26682 9417 26684
rect 9171 26630 9173 26682
rect 9353 26630 9355 26682
rect 9109 26628 9115 26630
rect 9171 26628 9195 26630
rect 9251 26628 9275 26630
rect 9331 26628 9355 26630
rect 9411 26628 9417 26630
rect 9109 26608 9417 26628
rect 8668 26580 8720 26586
rect 8668 26522 8720 26528
rect 8576 26036 8628 26042
rect 8576 25978 8628 25984
rect 9109 25596 9417 25616
rect 9109 25594 9115 25596
rect 9171 25594 9195 25596
rect 9251 25594 9275 25596
rect 9331 25594 9355 25596
rect 9411 25594 9417 25596
rect 9171 25542 9173 25594
rect 9353 25542 9355 25594
rect 9109 25540 9115 25542
rect 9171 25540 9195 25542
rect 9251 25540 9275 25542
rect 9331 25540 9355 25542
rect 9411 25540 9417 25542
rect 9109 25520 9417 25540
rect 9109 24508 9417 24528
rect 9109 24506 9115 24508
rect 9171 24506 9195 24508
rect 9251 24506 9275 24508
rect 9331 24506 9355 24508
rect 9411 24506 9417 24508
rect 9171 24454 9173 24506
rect 9353 24454 9355 24506
rect 9109 24452 9115 24454
rect 9171 24452 9195 24454
rect 9251 24452 9275 24454
rect 9331 24452 9355 24454
rect 9411 24452 9417 24454
rect 9109 24432 9417 24452
rect 9109 23420 9417 23440
rect 9109 23418 9115 23420
rect 9171 23418 9195 23420
rect 9251 23418 9275 23420
rect 9331 23418 9355 23420
rect 9411 23418 9417 23420
rect 9171 23366 9173 23418
rect 9353 23366 9355 23418
rect 9109 23364 9115 23366
rect 9171 23364 9195 23366
rect 9251 23364 9275 23366
rect 9331 23364 9355 23366
rect 9411 23364 9417 23366
rect 9109 23344 9417 23364
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 9140 22953 9168 23054
rect 9126 22944 9182 22953
rect 9126 22879 9182 22888
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 8864 22137 8892 22578
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 8850 22128 8906 22137
rect 8024 22092 8076 22098
rect 8850 22063 8906 22072
rect 8024 22034 8076 22040
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8956 21457 8984 21490
rect 8942 21448 8998 21457
rect 8942 21383 8998 21392
rect 9048 21026 9076 22374
rect 9109 22332 9417 22352
rect 9109 22330 9115 22332
rect 9171 22330 9195 22332
rect 9251 22330 9275 22332
rect 9331 22330 9355 22332
rect 9411 22330 9417 22332
rect 9171 22278 9173 22330
rect 9353 22278 9355 22330
rect 9109 22276 9115 22278
rect 9171 22276 9195 22278
rect 9251 22276 9275 22278
rect 9331 22276 9355 22278
rect 9411 22276 9417 22278
rect 9109 22256 9417 22276
rect 9508 22098 9536 42638
rect 9784 41614 9812 43590
rect 9876 42226 9904 44134
rect 9968 43314 9996 44678
rect 10140 44396 10192 44402
rect 10140 44338 10192 44344
rect 10152 44033 10180 44338
rect 10138 44024 10194 44033
rect 10138 43959 10194 43968
rect 10140 43784 10192 43790
rect 10140 43726 10192 43732
rect 10152 43353 10180 43726
rect 10138 43344 10194 43353
rect 9956 43308 10008 43314
rect 10138 43279 10194 43288
rect 9956 43250 10008 43256
rect 10140 42696 10192 42702
rect 10140 42638 10192 42644
rect 9956 42560 10008 42566
rect 10152 42537 10180 42638
rect 9956 42502 10008 42508
rect 10138 42528 10194 42537
rect 9864 42220 9916 42226
rect 9864 42162 9916 42168
rect 9864 42016 9916 42022
rect 9864 41958 9916 41964
rect 9772 41608 9824 41614
rect 9772 41550 9824 41556
rect 9876 40526 9904 41958
rect 9968 41138 9996 42502
rect 10138 42463 10194 42472
rect 10140 42220 10192 42226
rect 10140 42162 10192 42168
rect 10152 41857 10180 42162
rect 10138 41848 10194 41857
rect 10138 41783 10194 41792
rect 9956 41132 10008 41138
rect 9956 41074 10008 41080
rect 10140 41132 10192 41138
rect 10140 41074 10192 41080
rect 10152 41041 10180 41074
rect 10138 41032 10194 41041
rect 10138 40967 10194 40976
rect 9956 40928 10008 40934
rect 9956 40870 10008 40876
rect 9864 40520 9916 40526
rect 9864 40462 9916 40468
rect 9864 40384 9916 40390
rect 9864 40326 9916 40332
rect 9876 39438 9904 40326
rect 9968 40118 9996 40870
rect 10140 40520 10192 40526
rect 10140 40462 10192 40468
rect 10152 40361 10180 40462
rect 10138 40352 10194 40361
rect 10138 40287 10194 40296
rect 9956 40112 10008 40118
rect 9956 40054 10008 40060
rect 10140 40044 10192 40050
rect 10140 39986 10192 39992
rect 9956 39840 10008 39846
rect 9956 39782 10008 39788
rect 9864 39432 9916 39438
rect 9864 39374 9916 39380
rect 9864 38752 9916 38758
rect 9864 38694 9916 38700
rect 9876 37874 9904 38694
rect 9968 38350 9996 39782
rect 10152 39545 10180 39986
rect 10138 39536 10194 39545
rect 10138 39471 10194 39480
rect 10140 38956 10192 38962
rect 10140 38898 10192 38904
rect 10152 38729 10180 38898
rect 10138 38720 10194 38729
rect 10138 38655 10194 38664
rect 9956 38344 10008 38350
rect 9956 38286 10008 38292
rect 10140 38344 10192 38350
rect 10140 38286 10192 38292
rect 9956 38208 10008 38214
rect 9956 38150 10008 38156
rect 9864 37868 9916 37874
rect 9864 37810 9916 37816
rect 9968 37262 9996 38150
rect 10152 38049 10180 38286
rect 10138 38040 10194 38049
rect 10138 37975 10194 37984
rect 9956 37256 10008 37262
rect 10140 37256 10192 37262
rect 9956 37198 10008 37204
rect 10138 37224 10140 37233
rect 10192 37224 10194 37233
rect 10138 37159 10194 37168
rect 9956 37120 10008 37126
rect 9956 37062 10008 37068
rect 9968 36786 9996 37062
rect 9956 36780 10008 36786
rect 9956 36722 10008 36728
rect 10140 36780 10192 36786
rect 10140 36722 10192 36728
rect 10152 36553 10180 36722
rect 10138 36544 10194 36553
rect 10138 36479 10194 36488
rect 10140 36168 10192 36174
rect 10140 36110 10192 36116
rect 9956 36032 10008 36038
rect 9956 35974 10008 35980
rect 9968 35698 9996 35974
rect 10152 35737 10180 36110
rect 10138 35728 10194 35737
rect 9956 35692 10008 35698
rect 10138 35663 10194 35672
rect 9956 35634 10008 35640
rect 10140 35080 10192 35086
rect 10138 35048 10140 35057
rect 10192 35048 10194 35057
rect 10138 34983 10194 34992
rect 10140 34468 10192 34474
rect 10140 34410 10192 34416
rect 10152 34241 10180 34410
rect 10138 34232 10194 34241
rect 10138 34167 10194 34176
rect 10140 33992 10192 33998
rect 10140 33934 10192 33940
rect 9864 33856 9916 33862
rect 9864 33798 9916 33804
rect 9772 32224 9824 32230
rect 9772 32166 9824 32172
rect 9784 30734 9812 32166
rect 9876 31822 9904 33798
rect 10152 33561 10180 33934
rect 10138 33552 10194 33561
rect 10138 33487 10194 33496
rect 10140 32904 10192 32910
rect 10140 32846 10192 32852
rect 9956 32768 10008 32774
rect 10152 32745 10180 32846
rect 9956 32710 10008 32716
rect 10138 32736 10194 32745
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9968 31346 9996 32710
rect 10138 32671 10194 32680
rect 10140 32428 10192 32434
rect 10140 32370 10192 32376
rect 10152 31929 10180 32370
rect 10138 31920 10194 31929
rect 10138 31855 10194 31864
rect 9956 31340 10008 31346
rect 9956 31282 10008 31288
rect 10140 31340 10192 31346
rect 10140 31282 10192 31288
rect 10152 31249 10180 31282
rect 10138 31240 10194 31249
rect 10138 31175 10194 31184
rect 9864 31136 9916 31142
rect 9864 31078 9916 31084
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 9876 30258 9904 31078
rect 10140 30728 10192 30734
rect 10140 30670 10192 30676
rect 9956 30592 10008 30598
rect 9956 30534 10008 30540
rect 9864 30252 9916 30258
rect 9864 30194 9916 30200
rect 9864 30048 9916 30054
rect 9864 29990 9916 29996
rect 9680 29504 9732 29510
rect 9680 29446 9732 29452
rect 9692 29238 9720 29446
rect 9680 29232 9732 29238
rect 9680 29174 9732 29180
rect 9876 28966 9904 29990
rect 9968 29170 9996 30534
rect 10152 30433 10180 30670
rect 10138 30424 10194 30433
rect 10138 30359 10194 30368
rect 10140 30252 10192 30258
rect 10140 30194 10192 30200
rect 10152 29753 10180 30194
rect 10138 29744 10194 29753
rect 10138 29679 10194 29688
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 9956 29164 10008 29170
rect 9956 29106 10008 29112
rect 9956 29028 10008 29034
rect 9956 28970 10008 28976
rect 9864 28960 9916 28966
rect 9864 28902 9916 28908
rect 9968 28762 9996 28970
rect 10152 28937 10180 29582
rect 10138 28928 10194 28937
rect 10138 28863 10194 28872
rect 9956 28756 10008 28762
rect 9956 28698 10008 28704
rect 10140 28552 10192 28558
rect 10140 28494 10192 28500
rect 10152 28257 10180 28494
rect 10138 28248 10194 28257
rect 10138 28183 10194 28192
rect 10140 28076 10192 28082
rect 10140 28018 10192 28024
rect 9772 27872 9824 27878
rect 9772 27814 9824 27820
rect 9784 25974 9812 27814
rect 10152 27441 10180 28018
rect 10232 27464 10284 27470
rect 10138 27432 10194 27441
rect 10232 27406 10284 27412
rect 10138 27367 10194 27376
rect 9864 27328 9916 27334
rect 9864 27270 9916 27276
rect 9876 26586 9904 27270
rect 10048 26988 10100 26994
rect 10048 26930 10100 26936
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9864 26580 9916 26586
rect 9864 26522 9916 26528
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9876 25786 9904 26318
rect 9968 25974 9996 26726
rect 9956 25968 10008 25974
rect 10060 25945 10088 26930
rect 10244 26761 10272 27406
rect 10230 26752 10286 26761
rect 10230 26687 10286 26696
rect 10140 26444 10192 26450
rect 10140 26386 10192 26392
rect 10152 26042 10180 26386
rect 10140 26036 10192 26042
rect 10140 25978 10192 25984
rect 9956 25910 10008 25916
rect 10046 25936 10102 25945
rect 10046 25871 10102 25880
rect 9784 25758 9904 25786
rect 9784 25158 9812 25758
rect 10140 25288 10192 25294
rect 10138 25256 10140 25265
rect 10192 25256 10194 25265
rect 10138 25191 10194 25200
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 9784 23186 9812 25094
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 9876 23322 9904 24006
rect 9968 23730 9996 24550
rect 10152 24449 10180 24754
rect 10138 24440 10194 24449
rect 10138 24375 10194 24384
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 9956 23724 10008 23730
rect 9956 23666 10008 23672
rect 10152 23633 10180 24142
rect 10138 23624 10194 23633
rect 10138 23559 10194 23568
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9876 23066 9904 23258
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 9784 23038 9904 23066
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9496 22092 9548 22098
rect 9496 22034 9548 22040
rect 9600 21434 9628 22918
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9692 22030 9720 22714
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 9784 21554 9812 23038
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 9876 22030 9904 22918
rect 9968 22642 9996 22918
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 10060 22114 10088 23122
rect 10152 22642 10180 23462
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 9968 22086 10088 22114
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9772 21548 9824 21554
rect 9772 21490 9824 21496
rect 9876 21434 9904 21966
rect 9968 21570 9996 22086
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10060 21690 10088 21966
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 9968 21554 10088 21570
rect 9956 21548 10088 21554
rect 10008 21542 10088 21548
rect 9956 21490 10008 21496
rect 9600 21406 9720 21434
rect 9876 21406 9996 21434
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9109 21244 9417 21264
rect 9109 21242 9115 21244
rect 9171 21242 9195 21244
rect 9251 21242 9275 21244
rect 9331 21242 9355 21244
rect 9411 21242 9417 21244
rect 9171 21190 9173 21242
rect 9353 21190 9355 21242
rect 9109 21188 9115 21190
rect 9171 21188 9195 21190
rect 9251 21188 9275 21190
rect 9331 21188 9355 21190
rect 9411 21188 9417 21190
rect 9109 21168 9417 21188
rect 9048 20998 9168 21026
rect 9600 21010 9628 21286
rect 9036 20936 9088 20942
rect 9036 20878 9088 20884
rect 9048 20641 9076 20878
rect 9034 20632 9090 20641
rect 9034 20567 9090 20576
rect 9140 20534 9168 20998
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9692 20942 9720 21406
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9128 20528 9180 20534
rect 9128 20470 9180 20476
rect 9109 20156 9417 20176
rect 9109 20154 9115 20156
rect 9171 20154 9195 20156
rect 9251 20154 9275 20156
rect 9331 20154 9355 20156
rect 9411 20154 9417 20156
rect 9171 20102 9173 20154
rect 9353 20102 9355 20154
rect 9109 20100 9115 20102
rect 9171 20100 9195 20102
rect 9251 20100 9275 20102
rect 9331 20100 9355 20102
rect 9411 20100 9417 20102
rect 9109 20080 9417 20100
rect 9876 19514 9904 21286
rect 9968 21146 9996 21406
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 10060 20602 10088 21542
rect 10152 20942 10180 22578
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9968 20058 9996 20402
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 10138 19952 10194 19961
rect 10138 19887 10194 19896
rect 10152 19854 10180 19887
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 10244 19145 10272 19246
rect 10230 19136 10286 19145
rect 9109 19068 9417 19088
rect 10230 19071 10286 19080
rect 9109 19066 9115 19068
rect 9171 19066 9195 19068
rect 9251 19066 9275 19068
rect 9331 19066 9355 19068
rect 9411 19066 9417 19068
rect 9171 19014 9173 19066
rect 9353 19014 9355 19066
rect 9109 19012 9115 19014
rect 9171 19012 9195 19014
rect 9251 19012 9275 19014
rect 9331 19012 9355 19014
rect 9411 19012 9417 19014
rect 9109 18992 9417 19012
rect 9109 17980 9417 18000
rect 9109 17978 9115 17980
rect 9171 17978 9195 17980
rect 9251 17978 9275 17980
rect 9331 17978 9355 17980
rect 9411 17978 9417 17980
rect 9171 17926 9173 17978
rect 9353 17926 9355 17978
rect 9109 17924 9115 17926
rect 9171 17924 9195 17926
rect 9251 17924 9275 17926
rect 9331 17924 9355 17926
rect 9411 17924 9417 17926
rect 9109 17904 9417 17924
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7477 17436 7785 17456
rect 7477 17434 7483 17436
rect 7539 17434 7563 17436
rect 7619 17434 7643 17436
rect 7699 17434 7723 17436
rect 7779 17434 7785 17436
rect 7539 17382 7541 17434
rect 7721 17382 7723 17434
rect 7477 17380 7483 17382
rect 7539 17380 7563 17382
rect 7619 17380 7643 17382
rect 7699 17380 7723 17382
rect 7779 17380 7785 17382
rect 7477 17360 7785 17380
rect 9109 16892 9417 16912
rect 9109 16890 9115 16892
rect 9171 16890 9195 16892
rect 9251 16890 9275 16892
rect 9331 16890 9355 16892
rect 9411 16890 9417 16892
rect 9171 16838 9173 16890
rect 9353 16838 9355 16890
rect 9109 16836 9115 16838
rect 9171 16836 9195 16838
rect 9251 16836 9275 16838
rect 9331 16836 9355 16838
rect 9411 16836 9417 16838
rect 9109 16816 9417 16836
rect 7477 16348 7785 16368
rect 7477 16346 7483 16348
rect 7539 16346 7563 16348
rect 7619 16346 7643 16348
rect 7699 16346 7723 16348
rect 7779 16346 7785 16348
rect 7539 16294 7541 16346
rect 7721 16294 7723 16346
rect 7477 16292 7483 16294
rect 7539 16292 7563 16294
rect 7619 16292 7643 16294
rect 7699 16292 7723 16294
rect 7779 16292 7785 16294
rect 7477 16272 7785 16292
rect 9109 15804 9417 15824
rect 9109 15802 9115 15804
rect 9171 15802 9195 15804
rect 9251 15802 9275 15804
rect 9331 15802 9355 15804
rect 9411 15802 9417 15804
rect 9171 15750 9173 15802
rect 9353 15750 9355 15802
rect 9109 15748 9115 15750
rect 9171 15748 9195 15750
rect 9251 15748 9275 15750
rect 9331 15748 9355 15750
rect 9411 15748 9417 15750
rect 9109 15728 9417 15748
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 7477 15260 7785 15280
rect 7477 15258 7483 15260
rect 7539 15258 7563 15260
rect 7619 15258 7643 15260
rect 7699 15258 7723 15260
rect 7779 15258 7785 15260
rect 7539 15206 7541 15258
rect 7721 15206 7723 15258
rect 7477 15204 7483 15206
rect 7539 15204 7563 15206
rect 7619 15204 7643 15206
rect 7699 15204 7723 15206
rect 7779 15204 7785 15206
rect 7477 15184 7785 15204
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 5845 14716 6153 14736
rect 5845 14714 5851 14716
rect 5907 14714 5931 14716
rect 5987 14714 6011 14716
rect 6067 14714 6091 14716
rect 6147 14714 6153 14716
rect 5907 14662 5909 14714
rect 6089 14662 6091 14714
rect 5845 14660 5851 14662
rect 5907 14660 5931 14662
rect 5987 14660 6011 14662
rect 6067 14660 6091 14662
rect 6147 14660 6153 14662
rect 5845 14640 6153 14660
rect 9109 14716 9417 14736
rect 9109 14714 9115 14716
rect 9171 14714 9195 14716
rect 9251 14714 9275 14716
rect 9331 14714 9355 14716
rect 9411 14714 9417 14716
rect 9171 14662 9173 14714
rect 9353 14662 9355 14714
rect 9109 14660 9115 14662
rect 9171 14660 9195 14662
rect 9251 14660 9275 14662
rect 9331 14660 9355 14662
rect 9411 14660 9417 14662
rect 9109 14640 9417 14660
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 7477 14172 7785 14192
rect 7477 14170 7483 14172
rect 7539 14170 7563 14172
rect 7619 14170 7643 14172
rect 7699 14170 7723 14172
rect 7779 14170 7785 14172
rect 7539 14118 7541 14170
rect 7721 14118 7723 14170
rect 7477 14116 7483 14118
rect 7539 14116 7563 14118
rect 7619 14116 7643 14118
rect 7699 14116 7723 14118
rect 7779 14116 7785 14118
rect 7477 14096 7785 14116
rect 5845 13628 6153 13648
rect 5845 13626 5851 13628
rect 5907 13626 5931 13628
rect 5987 13626 6011 13628
rect 6067 13626 6091 13628
rect 6147 13626 6153 13628
rect 5907 13574 5909 13626
rect 6089 13574 6091 13626
rect 5845 13572 5851 13574
rect 5907 13572 5931 13574
rect 5987 13572 6011 13574
rect 6067 13572 6091 13574
rect 6147 13572 6153 13574
rect 5845 13552 6153 13572
rect 9109 13628 9417 13648
rect 9109 13626 9115 13628
rect 9171 13626 9195 13628
rect 9251 13626 9275 13628
rect 9331 13626 9355 13628
rect 9411 13626 9417 13628
rect 9171 13574 9173 13626
rect 9353 13574 9355 13626
rect 9109 13572 9115 13574
rect 9171 13572 9195 13574
rect 9251 13572 9275 13574
rect 9331 13572 9355 13574
rect 9411 13572 9417 13574
rect 9109 13552 9417 13572
rect 7477 13084 7785 13104
rect 7477 13082 7483 13084
rect 7539 13082 7563 13084
rect 7619 13082 7643 13084
rect 7699 13082 7723 13084
rect 7779 13082 7785 13084
rect 7539 13030 7541 13082
rect 7721 13030 7723 13082
rect 7477 13028 7483 13030
rect 7539 13028 7563 13030
rect 7619 13028 7643 13030
rect 7699 13028 7723 13030
rect 7779 13028 7785 13030
rect 7477 13008 7785 13028
rect 5845 12540 6153 12560
rect 5845 12538 5851 12540
rect 5907 12538 5931 12540
rect 5987 12538 6011 12540
rect 6067 12538 6091 12540
rect 6147 12538 6153 12540
rect 5907 12486 5909 12538
rect 6089 12486 6091 12538
rect 5845 12484 5851 12486
rect 5907 12484 5931 12486
rect 5987 12484 6011 12486
rect 6067 12484 6091 12486
rect 6147 12484 6153 12486
rect 5845 12464 6153 12484
rect 9109 12540 9417 12560
rect 9109 12538 9115 12540
rect 9171 12538 9195 12540
rect 9251 12538 9275 12540
rect 9331 12538 9355 12540
rect 9411 12538 9417 12540
rect 9171 12486 9173 12538
rect 9353 12486 9355 12538
rect 9109 12484 9115 12486
rect 9171 12484 9195 12486
rect 9251 12484 9275 12486
rect 9331 12484 9355 12486
rect 9411 12484 9417 12486
rect 9109 12464 9417 12484
rect 7477 11996 7785 12016
rect 7477 11994 7483 11996
rect 7539 11994 7563 11996
rect 7619 11994 7643 11996
rect 7699 11994 7723 11996
rect 7779 11994 7785 11996
rect 7539 11942 7541 11994
rect 7721 11942 7723 11994
rect 7477 11940 7483 11942
rect 7539 11940 7563 11942
rect 7619 11940 7643 11942
rect 7699 11940 7723 11942
rect 7779 11940 7785 11942
rect 7477 11920 7785 11940
rect 5845 11452 6153 11472
rect 5845 11450 5851 11452
rect 5907 11450 5931 11452
rect 5987 11450 6011 11452
rect 6067 11450 6091 11452
rect 6147 11450 6153 11452
rect 5907 11398 5909 11450
rect 6089 11398 6091 11450
rect 5845 11396 5851 11398
rect 5907 11396 5931 11398
rect 5987 11396 6011 11398
rect 6067 11396 6091 11398
rect 6147 11396 6153 11398
rect 5845 11376 6153 11396
rect 9109 11452 9417 11472
rect 9109 11450 9115 11452
rect 9171 11450 9195 11452
rect 9251 11450 9275 11452
rect 9331 11450 9355 11452
rect 9411 11450 9417 11452
rect 9171 11398 9173 11450
rect 9353 11398 9355 11450
rect 9109 11396 9115 11398
rect 9171 11396 9195 11398
rect 9251 11396 9275 11398
rect 9331 11396 9355 11398
rect 9411 11396 9417 11398
rect 9109 11376 9417 11396
rect 7477 10908 7785 10928
rect 7477 10906 7483 10908
rect 7539 10906 7563 10908
rect 7619 10906 7643 10908
rect 7699 10906 7723 10908
rect 7779 10906 7785 10908
rect 7539 10854 7541 10906
rect 7721 10854 7723 10906
rect 7477 10852 7483 10854
rect 7539 10852 7563 10854
rect 7619 10852 7643 10854
rect 7699 10852 7723 10854
rect 7779 10852 7785 10854
rect 7477 10832 7785 10852
rect 5845 10364 6153 10384
rect 5845 10362 5851 10364
rect 5907 10362 5931 10364
rect 5987 10362 6011 10364
rect 6067 10362 6091 10364
rect 6147 10362 6153 10364
rect 5907 10310 5909 10362
rect 6089 10310 6091 10362
rect 5845 10308 5851 10310
rect 5907 10308 5931 10310
rect 5987 10308 6011 10310
rect 6067 10308 6091 10310
rect 6147 10308 6153 10310
rect 5845 10288 6153 10308
rect 9109 10364 9417 10384
rect 9109 10362 9115 10364
rect 9171 10362 9195 10364
rect 9251 10362 9275 10364
rect 9331 10362 9355 10364
rect 9411 10362 9417 10364
rect 9171 10310 9173 10362
rect 9353 10310 9355 10362
rect 9109 10308 9115 10310
rect 9171 10308 9195 10310
rect 9251 10308 9275 10310
rect 9331 10308 9355 10310
rect 9411 10308 9417 10310
rect 9109 10288 9417 10308
rect 7477 9820 7785 9840
rect 7477 9818 7483 9820
rect 7539 9818 7563 9820
rect 7619 9818 7643 9820
rect 7699 9818 7723 9820
rect 7779 9818 7785 9820
rect 7539 9766 7541 9818
rect 7721 9766 7723 9818
rect 7477 9764 7483 9766
rect 7539 9764 7563 9766
rect 7619 9764 7643 9766
rect 7699 9764 7723 9766
rect 7779 9764 7785 9766
rect 7477 9744 7785 9764
rect 5845 9276 6153 9296
rect 5845 9274 5851 9276
rect 5907 9274 5931 9276
rect 5987 9274 6011 9276
rect 6067 9274 6091 9276
rect 6147 9274 6153 9276
rect 5907 9222 5909 9274
rect 6089 9222 6091 9274
rect 5845 9220 5851 9222
rect 5907 9220 5931 9222
rect 5987 9220 6011 9222
rect 6067 9220 6091 9222
rect 6147 9220 6153 9222
rect 5845 9200 6153 9220
rect 9109 9276 9417 9296
rect 9109 9274 9115 9276
rect 9171 9274 9195 9276
rect 9251 9274 9275 9276
rect 9331 9274 9355 9276
rect 9411 9274 9417 9276
rect 9171 9222 9173 9274
rect 9353 9222 9355 9274
rect 9109 9220 9115 9222
rect 9171 9220 9195 9222
rect 9251 9220 9275 9222
rect 9331 9220 9355 9222
rect 9411 9220 9417 9222
rect 9109 9200 9417 9220
rect 7477 8732 7785 8752
rect 7477 8730 7483 8732
rect 7539 8730 7563 8732
rect 7619 8730 7643 8732
rect 7699 8730 7723 8732
rect 7779 8730 7785 8732
rect 7539 8678 7541 8730
rect 7721 8678 7723 8730
rect 7477 8676 7483 8678
rect 7539 8676 7563 8678
rect 7619 8676 7643 8678
rect 7699 8676 7723 8678
rect 7779 8676 7785 8678
rect 7477 8656 7785 8676
rect 5845 8188 6153 8208
rect 5845 8186 5851 8188
rect 5907 8186 5931 8188
rect 5987 8186 6011 8188
rect 6067 8186 6091 8188
rect 6147 8186 6153 8188
rect 5907 8134 5909 8186
rect 6089 8134 6091 8186
rect 5845 8132 5851 8134
rect 5907 8132 5931 8134
rect 5987 8132 6011 8134
rect 6067 8132 6091 8134
rect 6147 8132 6153 8134
rect 5845 8112 6153 8132
rect 9109 8188 9417 8208
rect 9109 8186 9115 8188
rect 9171 8186 9195 8188
rect 9251 8186 9275 8188
rect 9331 8186 9355 8188
rect 9411 8186 9417 8188
rect 9171 8134 9173 8186
rect 9353 8134 9355 8186
rect 9109 8132 9115 8134
rect 9171 8132 9195 8134
rect 9251 8132 9275 8134
rect 9331 8132 9355 8134
rect 9411 8132 9417 8134
rect 9109 8112 9417 8132
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 7477 7644 7785 7664
rect 7477 7642 7483 7644
rect 7539 7642 7563 7644
rect 7619 7642 7643 7644
rect 7699 7642 7723 7644
rect 7779 7642 7785 7644
rect 7539 7590 7541 7642
rect 7721 7590 7723 7642
rect 7477 7588 7483 7590
rect 7539 7588 7563 7590
rect 7619 7588 7643 7590
rect 7699 7588 7723 7590
rect 7779 7588 7785 7590
rect 7477 7568 7785 7588
rect 5845 7100 6153 7120
rect 5845 7098 5851 7100
rect 5907 7098 5931 7100
rect 5987 7098 6011 7100
rect 6067 7098 6091 7100
rect 6147 7098 6153 7100
rect 5907 7046 5909 7098
rect 6089 7046 6091 7098
rect 5845 7044 5851 7046
rect 5907 7044 5931 7046
rect 5987 7044 6011 7046
rect 6067 7044 6091 7046
rect 6147 7044 6153 7046
rect 5845 7024 6153 7044
rect 9109 7100 9417 7120
rect 9109 7098 9115 7100
rect 9171 7098 9195 7100
rect 9251 7098 9275 7100
rect 9331 7098 9355 7100
rect 9411 7098 9417 7100
rect 9171 7046 9173 7098
rect 9353 7046 9355 7098
rect 9109 7044 9115 7046
rect 9171 7044 9195 7046
rect 9251 7044 9275 7046
rect 9331 7044 9355 7046
rect 9411 7044 9417 7046
rect 9109 7024 9417 7044
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 7477 6556 7785 6576
rect 7477 6554 7483 6556
rect 7539 6554 7563 6556
rect 7619 6554 7643 6556
rect 7699 6554 7723 6556
rect 7779 6554 7785 6556
rect 7539 6502 7541 6554
rect 7721 6502 7723 6554
rect 7477 6500 7483 6502
rect 7539 6500 7563 6502
rect 7619 6500 7643 6502
rect 7699 6500 7723 6502
rect 7779 6500 7785 6502
rect 7477 6480 7785 6500
rect 9968 6390 9996 6598
rect 9956 6384 10008 6390
rect 10152 6361 10180 6734
rect 9956 6326 10008 6332
rect 10138 6352 10194 6361
rect 10138 6287 10194 6296
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 5845 6012 6153 6032
rect 5845 6010 5851 6012
rect 5907 6010 5931 6012
rect 5987 6010 6011 6012
rect 6067 6010 6091 6012
rect 6147 6010 6153 6012
rect 5907 5958 5909 6010
rect 6089 5958 6091 6010
rect 5845 5956 5851 5958
rect 5907 5956 5931 5958
rect 5987 5956 6011 5958
rect 6067 5956 6091 5958
rect 6147 5956 6153 5958
rect 5845 5936 6153 5956
rect 9109 6012 9417 6032
rect 9109 6010 9115 6012
rect 9171 6010 9195 6012
rect 9251 6010 9275 6012
rect 9331 6010 9355 6012
rect 9411 6010 9417 6012
rect 9171 5958 9173 6010
rect 9353 5958 9355 6010
rect 9109 5956 9115 5958
rect 9171 5956 9195 5958
rect 9251 5956 9275 5958
rect 9331 5956 9355 5958
rect 9411 5956 9417 5958
rect 9109 5936 9417 5956
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4213 5468 4521 5488
rect 4213 5466 4219 5468
rect 4275 5466 4299 5468
rect 4355 5466 4379 5468
rect 4435 5466 4459 5468
rect 4515 5466 4521 5468
rect 4275 5414 4277 5466
rect 4457 5414 4459 5466
rect 4213 5412 4219 5414
rect 4275 5412 4299 5414
rect 4355 5412 4379 5414
rect 4435 5412 4459 5414
rect 4515 5412 4521 5414
rect 4213 5392 4521 5412
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 4080 4282 4108 5170
rect 4632 4622 4660 5850
rect 4724 5166 4752 5850
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 7477 5468 7785 5488
rect 7477 5466 7483 5468
rect 7539 5466 7563 5468
rect 7619 5466 7643 5468
rect 7699 5466 7723 5468
rect 7779 5466 7785 5468
rect 7539 5414 7541 5466
rect 7721 5414 7723 5466
rect 7477 5412 7483 5414
rect 7539 5412 7563 5414
rect 7619 5412 7643 5414
rect 7699 5412 7723 5414
rect 7779 5412 7785 5414
rect 7477 5392 7785 5412
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 5845 4924 6153 4944
rect 5845 4922 5851 4924
rect 5907 4922 5931 4924
rect 5987 4922 6011 4924
rect 6067 4922 6091 4924
rect 6147 4922 6153 4924
rect 5907 4870 5909 4922
rect 6089 4870 6091 4922
rect 5845 4868 5851 4870
rect 5907 4868 5931 4870
rect 5987 4868 6011 4870
rect 6067 4868 6091 4870
rect 6147 4868 6153 4870
rect 5845 4848 6153 4868
rect 9109 4924 9417 4944
rect 9109 4922 9115 4924
rect 9171 4922 9195 4924
rect 9251 4922 9275 4924
rect 9331 4922 9355 4924
rect 9411 4922 9417 4924
rect 9171 4870 9173 4922
rect 9353 4870 9355 4922
rect 9109 4868 9115 4870
rect 9171 4868 9195 4870
rect 9251 4868 9275 4870
rect 9331 4868 9355 4870
rect 9411 4868 9417 4870
rect 9109 4848 9417 4868
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4213 4380 4521 4400
rect 4213 4378 4219 4380
rect 4275 4378 4299 4380
rect 4355 4378 4379 4380
rect 4435 4378 4459 4380
rect 4515 4378 4521 4380
rect 4275 4326 4277 4378
rect 4457 4326 4459 4378
rect 4213 4324 4219 4326
rect 4275 4324 4299 4326
rect 4355 4324 4379 4326
rect 4435 4324 4459 4326
rect 4515 4324 4521 4326
rect 4213 4304 4521 4324
rect 7477 4380 7785 4400
rect 7477 4378 7483 4380
rect 7539 4378 7563 4380
rect 7619 4378 7643 4380
rect 7699 4378 7723 4380
rect 7779 4378 7785 4380
rect 7539 4326 7541 4378
rect 7721 4326 7723 4378
rect 7477 4324 7483 4326
rect 7539 4324 7563 4326
rect 7619 4324 7643 4326
rect 7699 4324 7723 4326
rect 7779 4324 7785 4326
rect 7477 4304 7785 4324
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 5845 3836 6153 3856
rect 5845 3834 5851 3836
rect 5907 3834 5931 3836
rect 5987 3834 6011 3836
rect 6067 3834 6091 3836
rect 6147 3834 6153 3836
rect 5907 3782 5909 3834
rect 6089 3782 6091 3834
rect 5845 3780 5851 3782
rect 5907 3780 5931 3782
rect 5987 3780 6011 3782
rect 6067 3780 6091 3782
rect 6147 3780 6153 3782
rect 5845 3760 6153 3780
rect 9109 3836 9417 3856
rect 9109 3834 9115 3836
rect 9171 3834 9195 3836
rect 9251 3834 9275 3836
rect 9331 3834 9355 3836
rect 9411 3834 9417 3836
rect 9171 3782 9173 3834
rect 9353 3782 9355 3834
rect 9109 3780 9115 3782
rect 9171 3780 9195 3782
rect 9251 3780 9275 3782
rect 9331 3780 9355 3782
rect 9411 3780 9417 3782
rect 9109 3760 9417 3780
rect 9876 3738 9904 5646
rect 9968 5370 9996 6190
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10152 5545 10180 5646
rect 10138 5536 10194 5545
rect 10138 5471 10194 5480
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10152 4865 10180 5170
rect 10138 4856 10194 4865
rect 10138 4791 10194 4800
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10152 4049 10180 4082
rect 10138 4040 10194 4049
rect 10138 3975 10194 3984
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 4213 3292 4521 3312
rect 4213 3290 4219 3292
rect 4275 3290 4299 3292
rect 4355 3290 4379 3292
rect 4435 3290 4459 3292
rect 4515 3290 4521 3292
rect 4275 3238 4277 3290
rect 4457 3238 4459 3290
rect 4213 3236 4219 3238
rect 4275 3236 4299 3238
rect 4355 3236 4379 3238
rect 4435 3236 4459 3238
rect 4515 3236 4521 3238
rect 4213 3216 4521 3236
rect 7477 3292 7785 3312
rect 7477 3290 7483 3292
rect 7539 3290 7563 3292
rect 7619 3290 7643 3292
rect 7699 3290 7723 3292
rect 7779 3290 7785 3292
rect 7539 3238 7541 3290
rect 7721 3238 7723 3290
rect 7477 3236 7483 3238
rect 7539 3236 7563 3238
rect 7619 3236 7643 3238
rect 7699 3236 7723 3238
rect 7779 3236 7785 3238
rect 7477 3216 7785 3236
rect 9876 3058 9904 3470
rect 10152 3369 10180 3470
rect 10138 3360 10194 3369
rect 10138 3295 10194 3304
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 2582 2748 2890 2768
rect 2582 2746 2588 2748
rect 2644 2746 2668 2748
rect 2724 2746 2748 2748
rect 2804 2746 2828 2748
rect 2884 2746 2890 2748
rect 2644 2694 2646 2746
rect 2826 2694 2828 2746
rect 2582 2692 2588 2694
rect 2644 2692 2668 2694
rect 2724 2692 2748 2694
rect 2804 2692 2828 2694
rect 2884 2692 2890 2694
rect 2582 2672 2890 2692
rect 2976 2746 3188 2774
rect 5845 2748 6153 2768
rect 5845 2746 5851 2748
rect 5907 2746 5931 2748
rect 5987 2746 6011 2748
rect 6067 2746 6091 2748
rect 6147 2746 6153 2748
rect 2976 2446 3004 2746
rect 5907 2694 5909 2746
rect 6089 2694 6091 2746
rect 5845 2692 5851 2694
rect 5907 2692 5931 2694
rect 5987 2692 6011 2694
rect 6067 2692 6091 2694
rect 6147 2692 6153 2694
rect 5845 2672 6153 2692
rect 9109 2748 9417 2768
rect 9109 2746 9115 2748
rect 9171 2746 9195 2748
rect 9251 2746 9275 2748
rect 9331 2746 9355 2748
rect 9411 2746 9417 2748
rect 9171 2694 9173 2746
rect 9353 2694 9355 2746
rect 9109 2692 9115 2694
rect 9171 2692 9195 2694
rect 9251 2692 9275 2694
rect 9331 2692 9355 2694
rect 9411 2692 9417 2694
rect 9109 2672 9417 2692
rect 10152 2553 10180 2926
rect 10138 2544 10194 2553
rect 10138 2479 10194 2488
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 1490 2000 1546 2009
rect 1490 1935 1546 1944
rect 1398 912 1454 921
rect 1398 847 1454 856
rect 2792 377 2820 2246
rect 3068 1465 3096 2246
rect 4213 2204 4521 2224
rect 4213 2202 4219 2204
rect 4275 2202 4299 2204
rect 4355 2202 4379 2204
rect 4435 2202 4459 2204
rect 4515 2202 4521 2204
rect 4275 2150 4277 2202
rect 4457 2150 4459 2202
rect 4213 2148 4219 2150
rect 4275 2148 4299 2150
rect 4355 2148 4379 2150
rect 4435 2148 4459 2150
rect 4515 2148 4521 2150
rect 4213 2128 4521 2148
rect 7477 2204 7785 2224
rect 7477 2202 7483 2204
rect 7539 2202 7563 2204
rect 7619 2202 7643 2204
rect 7699 2202 7723 2204
rect 7779 2202 7785 2204
rect 7539 2150 7541 2202
rect 7721 2150 7723 2202
rect 7477 2148 7483 2150
rect 7539 2148 7563 2150
rect 7619 2148 7643 2150
rect 7699 2148 7723 2150
rect 7779 2148 7785 2150
rect 7477 2128 7785 2148
rect 10152 1873 10180 2382
rect 10138 1864 10194 1873
rect 10138 1799 10194 1808
rect 3054 1456 3110 1465
rect 3054 1391 3110 1400
rect 2778 368 2834 377
rect 2778 303 2834 312
<< via2 >>
rect 3790 79600 3846 79656
rect 3054 79056 3110 79112
rect 1490 78512 1546 78568
rect 2962 77968 3018 78024
rect 2588 77818 2644 77820
rect 2668 77818 2724 77820
rect 2748 77818 2804 77820
rect 2828 77818 2884 77820
rect 2588 77766 2634 77818
rect 2634 77766 2644 77818
rect 2668 77766 2698 77818
rect 2698 77766 2710 77818
rect 2710 77766 2724 77818
rect 2748 77766 2762 77818
rect 2762 77766 2774 77818
rect 2774 77766 2804 77818
rect 2828 77766 2838 77818
rect 2838 77766 2884 77818
rect 2588 77764 2644 77766
rect 2668 77764 2724 77766
rect 2748 77764 2804 77766
rect 2828 77764 2884 77766
rect 1398 76880 1454 76936
rect 1306 76336 1362 76392
rect 1398 75792 1454 75848
rect 1306 74704 1362 74760
rect 1398 73616 1454 73672
rect 2042 77460 2044 77480
rect 2044 77460 2096 77480
rect 2096 77460 2098 77480
rect 2042 77424 2098 77460
rect 2042 75284 2044 75304
rect 2044 75284 2096 75304
rect 2096 75284 2098 75304
rect 2042 75248 2098 75284
rect 9586 79464 9642 79520
rect 9494 77968 9550 78024
rect 5851 77818 5907 77820
rect 5931 77818 5987 77820
rect 6011 77818 6067 77820
rect 6091 77818 6147 77820
rect 5851 77766 5897 77818
rect 5897 77766 5907 77818
rect 5931 77766 5961 77818
rect 5961 77766 5973 77818
rect 5973 77766 5987 77818
rect 6011 77766 6025 77818
rect 6025 77766 6037 77818
rect 6037 77766 6067 77818
rect 6091 77766 6101 77818
rect 6101 77766 6147 77818
rect 5851 77764 5907 77766
rect 5931 77764 5987 77766
rect 6011 77764 6067 77766
rect 6091 77764 6147 77766
rect 9115 77818 9171 77820
rect 9195 77818 9251 77820
rect 9275 77818 9331 77820
rect 9355 77818 9411 77820
rect 9115 77766 9161 77818
rect 9161 77766 9171 77818
rect 9195 77766 9225 77818
rect 9225 77766 9237 77818
rect 9237 77766 9251 77818
rect 9275 77766 9289 77818
rect 9289 77766 9301 77818
rect 9301 77766 9331 77818
rect 9355 77766 9365 77818
rect 9365 77766 9411 77818
rect 9115 77764 9171 77766
rect 9195 77764 9251 77766
rect 9275 77764 9331 77766
rect 9355 77764 9411 77766
rect 2588 76730 2644 76732
rect 2668 76730 2724 76732
rect 2748 76730 2804 76732
rect 2828 76730 2884 76732
rect 2588 76678 2634 76730
rect 2634 76678 2644 76730
rect 2668 76678 2698 76730
rect 2698 76678 2710 76730
rect 2710 76678 2724 76730
rect 2748 76678 2762 76730
rect 2762 76678 2774 76730
rect 2774 76678 2804 76730
rect 2828 76678 2838 76730
rect 2838 76678 2884 76730
rect 2588 76676 2644 76678
rect 2668 76676 2724 76678
rect 2748 76676 2804 76678
rect 2828 76676 2884 76678
rect 2588 75642 2644 75644
rect 2668 75642 2724 75644
rect 2748 75642 2804 75644
rect 2828 75642 2884 75644
rect 2588 75590 2634 75642
rect 2634 75590 2644 75642
rect 2668 75590 2698 75642
rect 2698 75590 2710 75642
rect 2710 75590 2724 75642
rect 2748 75590 2762 75642
rect 2762 75590 2774 75642
rect 2774 75590 2804 75642
rect 2828 75590 2838 75642
rect 2838 75590 2884 75642
rect 2588 75588 2644 75590
rect 2668 75588 2724 75590
rect 2748 75588 2804 75590
rect 2828 75588 2884 75590
rect 2588 74554 2644 74556
rect 2668 74554 2724 74556
rect 2748 74554 2804 74556
rect 2828 74554 2884 74556
rect 2588 74502 2634 74554
rect 2634 74502 2644 74554
rect 2668 74502 2698 74554
rect 2698 74502 2710 74554
rect 2710 74502 2724 74554
rect 2748 74502 2762 74554
rect 2762 74502 2774 74554
rect 2774 74502 2804 74554
rect 2828 74502 2838 74554
rect 2838 74502 2884 74554
rect 2588 74500 2644 74502
rect 2668 74500 2724 74502
rect 2748 74500 2804 74502
rect 2828 74500 2884 74502
rect 2588 73466 2644 73468
rect 2668 73466 2724 73468
rect 2748 73466 2804 73468
rect 2828 73466 2884 73468
rect 2588 73414 2634 73466
rect 2634 73414 2644 73466
rect 2668 73414 2698 73466
rect 2698 73414 2710 73466
rect 2710 73414 2724 73466
rect 2748 73414 2762 73466
rect 2762 73414 2774 73466
rect 2774 73414 2804 73466
rect 2828 73414 2838 73466
rect 2838 73414 2884 73466
rect 2588 73412 2644 73414
rect 2668 73412 2724 73414
rect 2748 73412 2804 73414
rect 2828 73412 2884 73414
rect 2042 72936 2098 72992
rect 1398 72392 1454 72448
rect 1398 71848 1454 71904
rect 1398 71304 1454 71360
rect 1398 70760 1454 70816
rect 1398 70216 1454 70272
rect 1398 69672 1454 69728
rect 1398 69128 1454 69184
rect 1398 68584 1454 68640
rect 1398 68040 1454 68096
rect 1214 65728 1270 65784
rect 1398 66272 1454 66328
rect 1306 65184 1362 65240
rect 1398 64640 1454 64696
rect 1490 63980 1546 64016
rect 1490 63960 1492 63980
rect 1492 63960 1544 63980
rect 1544 63960 1546 63980
rect 1306 63552 1362 63608
rect 1490 61376 1546 61432
rect 1398 60832 1454 60888
rect 1490 60288 1546 60344
rect 1398 59608 1454 59664
rect 1490 59064 1546 59120
rect 1398 58520 1454 58576
rect 1490 57976 1546 58032
rect 2588 72378 2644 72380
rect 2668 72378 2724 72380
rect 2748 72378 2804 72380
rect 2828 72378 2884 72380
rect 2588 72326 2634 72378
rect 2634 72326 2644 72378
rect 2668 72326 2698 72378
rect 2698 72326 2710 72378
rect 2710 72326 2724 72378
rect 2748 72326 2762 72378
rect 2762 72326 2774 72378
rect 2774 72326 2804 72378
rect 2828 72326 2838 72378
rect 2838 72326 2884 72378
rect 2588 72324 2644 72326
rect 2668 72324 2724 72326
rect 2748 72324 2804 72326
rect 2828 72324 2884 72326
rect 1582 57704 1638 57760
rect 1398 56888 1454 56944
rect 1490 54168 1546 54224
rect 1490 53624 1546 53680
rect 1490 52944 1546 53000
rect 1490 52400 1546 52456
rect 1490 51312 1546 51368
rect 1674 50940 1676 50960
rect 1676 50940 1728 50960
rect 1728 50940 1730 50960
rect 1674 50904 1730 50940
rect 2226 67496 2282 67552
rect 2226 66952 2282 67008
rect 2588 71290 2644 71292
rect 2668 71290 2724 71292
rect 2748 71290 2804 71292
rect 2828 71290 2884 71292
rect 2588 71238 2634 71290
rect 2634 71238 2644 71290
rect 2668 71238 2698 71290
rect 2698 71238 2710 71290
rect 2710 71238 2724 71290
rect 2748 71238 2762 71290
rect 2762 71238 2774 71290
rect 2774 71238 2804 71290
rect 2828 71238 2838 71290
rect 2838 71238 2884 71290
rect 2588 71236 2644 71238
rect 2668 71236 2724 71238
rect 2748 71236 2804 71238
rect 2828 71236 2884 71238
rect 2588 70202 2644 70204
rect 2668 70202 2724 70204
rect 2748 70202 2804 70204
rect 2828 70202 2884 70204
rect 2588 70150 2634 70202
rect 2634 70150 2644 70202
rect 2668 70150 2698 70202
rect 2698 70150 2710 70202
rect 2710 70150 2724 70202
rect 2748 70150 2762 70202
rect 2762 70150 2774 70202
rect 2774 70150 2804 70202
rect 2828 70150 2838 70202
rect 2838 70150 2884 70202
rect 2588 70148 2644 70150
rect 2668 70148 2724 70150
rect 2748 70148 2804 70150
rect 2828 70148 2884 70150
rect 2588 69114 2644 69116
rect 2668 69114 2724 69116
rect 2748 69114 2804 69116
rect 2828 69114 2884 69116
rect 2588 69062 2634 69114
rect 2634 69062 2644 69114
rect 2668 69062 2698 69114
rect 2698 69062 2710 69114
rect 2710 69062 2724 69114
rect 2748 69062 2762 69114
rect 2762 69062 2774 69114
rect 2774 69062 2804 69114
rect 2828 69062 2838 69114
rect 2838 69062 2884 69114
rect 2588 69060 2644 69062
rect 2668 69060 2724 69062
rect 2748 69060 2804 69062
rect 2828 69060 2884 69062
rect 4219 77274 4275 77276
rect 4299 77274 4355 77276
rect 4379 77274 4435 77276
rect 4459 77274 4515 77276
rect 4219 77222 4265 77274
rect 4265 77222 4275 77274
rect 4299 77222 4329 77274
rect 4329 77222 4341 77274
rect 4341 77222 4355 77274
rect 4379 77222 4393 77274
rect 4393 77222 4405 77274
rect 4405 77222 4435 77274
rect 4459 77222 4469 77274
rect 4469 77222 4515 77274
rect 4219 77220 4275 77222
rect 4299 77220 4355 77222
rect 4379 77220 4435 77222
rect 4459 77220 4515 77222
rect 4219 76186 4275 76188
rect 4299 76186 4355 76188
rect 4379 76186 4435 76188
rect 4459 76186 4515 76188
rect 4219 76134 4265 76186
rect 4265 76134 4275 76186
rect 4299 76134 4329 76186
rect 4329 76134 4341 76186
rect 4341 76134 4355 76186
rect 4379 76134 4393 76186
rect 4393 76134 4405 76186
rect 4405 76134 4435 76186
rect 4459 76134 4469 76186
rect 4469 76134 4515 76186
rect 4219 76132 4275 76134
rect 4299 76132 4355 76134
rect 4379 76132 4435 76134
rect 4459 76132 4515 76134
rect 4219 75098 4275 75100
rect 4299 75098 4355 75100
rect 4379 75098 4435 75100
rect 4459 75098 4515 75100
rect 4219 75046 4265 75098
rect 4265 75046 4275 75098
rect 4299 75046 4329 75098
rect 4329 75046 4341 75098
rect 4341 75046 4355 75098
rect 4379 75046 4393 75098
rect 4393 75046 4405 75098
rect 4405 75046 4435 75098
rect 4459 75046 4469 75098
rect 4469 75046 4515 75098
rect 4219 75044 4275 75046
rect 4299 75044 4355 75046
rect 4379 75044 4435 75046
rect 4459 75044 4515 75046
rect 7483 77274 7539 77276
rect 7563 77274 7619 77276
rect 7643 77274 7699 77276
rect 7723 77274 7779 77276
rect 7483 77222 7529 77274
rect 7529 77222 7539 77274
rect 7563 77222 7593 77274
rect 7593 77222 7605 77274
rect 7605 77222 7619 77274
rect 7643 77222 7657 77274
rect 7657 77222 7669 77274
rect 7669 77222 7699 77274
rect 7723 77222 7733 77274
rect 7733 77222 7779 77274
rect 7483 77220 7539 77222
rect 7563 77220 7619 77222
rect 7643 77220 7699 77222
rect 7723 77220 7779 77222
rect 10966 78668 11022 78704
rect 10966 78648 10968 78668
rect 10968 78648 11020 78668
rect 11020 78648 11022 78668
rect 10046 77152 10102 77208
rect 5851 76730 5907 76732
rect 5931 76730 5987 76732
rect 6011 76730 6067 76732
rect 6091 76730 6147 76732
rect 5851 76678 5897 76730
rect 5897 76678 5907 76730
rect 5931 76678 5961 76730
rect 5961 76678 5973 76730
rect 5973 76678 5987 76730
rect 6011 76678 6025 76730
rect 6025 76678 6037 76730
rect 6037 76678 6067 76730
rect 6091 76678 6101 76730
rect 6101 76678 6147 76730
rect 5851 76676 5907 76678
rect 5931 76676 5987 76678
rect 6011 76676 6067 76678
rect 6091 76676 6147 76678
rect 7483 76186 7539 76188
rect 7563 76186 7619 76188
rect 7643 76186 7699 76188
rect 7723 76186 7779 76188
rect 7483 76134 7529 76186
rect 7529 76134 7539 76186
rect 7563 76134 7593 76186
rect 7593 76134 7605 76186
rect 7605 76134 7619 76186
rect 7643 76134 7657 76186
rect 7657 76134 7669 76186
rect 7669 76134 7699 76186
rect 7723 76134 7733 76186
rect 7733 76134 7779 76186
rect 7483 76132 7539 76134
rect 7563 76132 7619 76134
rect 7643 76132 7699 76134
rect 7723 76132 7779 76134
rect 5851 75642 5907 75644
rect 5931 75642 5987 75644
rect 6011 75642 6067 75644
rect 6091 75642 6147 75644
rect 5851 75590 5897 75642
rect 5897 75590 5907 75642
rect 5931 75590 5961 75642
rect 5961 75590 5973 75642
rect 5973 75590 5987 75642
rect 6011 75590 6025 75642
rect 6025 75590 6037 75642
rect 6037 75590 6067 75642
rect 6091 75590 6101 75642
rect 6101 75590 6147 75642
rect 5851 75588 5907 75590
rect 5931 75588 5987 75590
rect 6011 75588 6067 75590
rect 6091 75588 6147 75590
rect 7483 75098 7539 75100
rect 7563 75098 7619 75100
rect 7643 75098 7699 75100
rect 7723 75098 7779 75100
rect 7483 75046 7529 75098
rect 7529 75046 7539 75098
rect 7563 75046 7593 75098
rect 7593 75046 7605 75098
rect 7605 75046 7619 75098
rect 7643 75046 7657 75098
rect 7657 75046 7669 75098
rect 7669 75046 7699 75098
rect 7723 75046 7733 75098
rect 7733 75046 7779 75098
rect 7483 75044 7539 75046
rect 7563 75044 7619 75046
rect 7643 75044 7699 75046
rect 7723 75044 7779 75046
rect 5851 74554 5907 74556
rect 5931 74554 5987 74556
rect 6011 74554 6067 74556
rect 6091 74554 6147 74556
rect 5851 74502 5897 74554
rect 5897 74502 5907 74554
rect 5931 74502 5961 74554
rect 5961 74502 5973 74554
rect 5973 74502 5987 74554
rect 6011 74502 6025 74554
rect 6025 74502 6037 74554
rect 6037 74502 6067 74554
rect 6091 74502 6101 74554
rect 6101 74502 6147 74554
rect 5851 74500 5907 74502
rect 5931 74500 5987 74502
rect 6011 74500 6067 74502
rect 6091 74500 6147 74502
rect 3790 74196 3792 74216
rect 3792 74196 3844 74216
rect 3844 74196 3846 74216
rect 3790 74160 3846 74196
rect 2588 68026 2644 68028
rect 2668 68026 2724 68028
rect 2748 68026 2804 68028
rect 2828 68026 2884 68028
rect 2588 67974 2634 68026
rect 2634 67974 2644 68026
rect 2668 67974 2698 68026
rect 2698 67974 2710 68026
rect 2710 67974 2724 68026
rect 2748 67974 2762 68026
rect 2762 67974 2774 68026
rect 2774 67974 2804 68026
rect 2828 67974 2838 68026
rect 2838 67974 2884 68026
rect 2588 67972 2644 67974
rect 2668 67972 2724 67974
rect 2748 67972 2804 67974
rect 2828 67972 2884 67974
rect 2588 66938 2644 66940
rect 2668 66938 2724 66940
rect 2748 66938 2804 66940
rect 2828 66938 2884 66940
rect 2588 66886 2634 66938
rect 2634 66886 2644 66938
rect 2668 66886 2698 66938
rect 2698 66886 2710 66938
rect 2710 66886 2724 66938
rect 2748 66886 2762 66938
rect 2762 66886 2774 66938
rect 2774 66886 2804 66938
rect 2828 66886 2838 66938
rect 2838 66886 2884 66938
rect 2588 66884 2644 66886
rect 2668 66884 2724 66886
rect 2748 66884 2804 66886
rect 2828 66884 2884 66886
rect 1950 57840 2006 57896
rect 2588 65850 2644 65852
rect 2668 65850 2724 65852
rect 2748 65850 2804 65852
rect 2828 65850 2884 65852
rect 2588 65798 2634 65850
rect 2634 65798 2644 65850
rect 2668 65798 2698 65850
rect 2698 65798 2710 65850
rect 2710 65798 2724 65850
rect 2748 65798 2762 65850
rect 2762 65798 2774 65850
rect 2774 65798 2804 65850
rect 2828 65798 2838 65850
rect 2838 65798 2884 65850
rect 2588 65796 2644 65798
rect 2668 65796 2724 65798
rect 2748 65796 2804 65798
rect 2828 65796 2884 65798
rect 2588 64762 2644 64764
rect 2668 64762 2724 64764
rect 2748 64762 2804 64764
rect 2828 64762 2884 64764
rect 2588 64710 2634 64762
rect 2634 64710 2644 64762
rect 2668 64710 2698 64762
rect 2698 64710 2710 64762
rect 2710 64710 2724 64762
rect 2748 64710 2762 64762
rect 2762 64710 2774 64762
rect 2774 64710 2804 64762
rect 2828 64710 2838 64762
rect 2838 64710 2884 64762
rect 2588 64708 2644 64710
rect 2668 64708 2724 64710
rect 2748 64708 2804 64710
rect 2828 64708 2884 64710
rect 2778 64096 2834 64152
rect 2502 63980 2558 64016
rect 2502 63960 2504 63980
rect 2504 63960 2556 63980
rect 2556 63960 2558 63980
rect 2588 63674 2644 63676
rect 2668 63674 2724 63676
rect 2748 63674 2804 63676
rect 2828 63674 2884 63676
rect 2588 63622 2634 63674
rect 2634 63622 2644 63674
rect 2668 63622 2698 63674
rect 2698 63622 2710 63674
rect 2710 63622 2724 63674
rect 2748 63622 2762 63674
rect 2762 63622 2774 63674
rect 2774 63622 2804 63674
rect 2828 63622 2838 63674
rect 2838 63622 2884 63674
rect 2588 63620 2644 63622
rect 2668 63620 2724 63622
rect 2748 63620 2804 63622
rect 2828 63620 2884 63622
rect 2318 61920 2374 61976
rect 2226 59336 2282 59392
rect 1490 49700 1546 49736
rect 1490 49680 1492 49700
rect 1492 49680 1544 49700
rect 1544 49680 1546 49700
rect 1490 49136 1546 49192
rect 1490 48612 1546 48648
rect 1490 48592 1492 48612
rect 1492 48592 1544 48612
rect 1544 48592 1546 48612
rect 1490 48048 1546 48104
rect 1490 47524 1546 47560
rect 1490 47504 1492 47524
rect 1492 47504 1544 47524
rect 1544 47504 1546 47524
rect 1490 46960 1546 47016
rect 1490 46316 1492 46336
rect 1492 46316 1544 46336
rect 1544 46316 1546 46336
rect 1490 46280 1546 46316
rect 1490 45772 1492 45792
rect 1492 45772 1544 45792
rect 1544 45772 1546 45792
rect 1490 45736 1546 45772
rect 1490 45228 1492 45248
rect 1492 45228 1544 45248
rect 1544 45228 1546 45248
rect 1490 45192 1546 45228
rect 1490 44684 1492 44704
rect 1492 44684 1544 44704
rect 1544 44684 1546 44704
rect 1490 44648 1546 44684
rect 1490 44140 1492 44160
rect 1492 44140 1544 44160
rect 1544 44140 1546 44160
rect 1490 44104 1546 44140
rect 1490 43596 1492 43616
rect 1492 43596 1544 43616
rect 1544 43596 1546 43616
rect 1490 43560 1546 43596
rect 1490 43052 1492 43072
rect 1492 43052 1544 43072
rect 1544 43052 1546 43072
rect 1490 43016 1546 43052
rect 1490 42508 1492 42528
rect 1492 42508 1544 42528
rect 1544 42508 1546 42528
rect 1490 42472 1546 42508
rect 1490 41964 1492 41984
rect 1492 41964 1544 41984
rect 1544 41964 1546 41984
rect 1490 41928 1546 41964
rect 1490 41420 1492 41440
rect 1492 41420 1544 41440
rect 1544 41420 1546 41440
rect 1490 41384 1546 41420
rect 1490 40876 1492 40896
rect 1492 40876 1544 40896
rect 1544 40876 1546 40896
rect 1490 40840 1546 40876
rect 1490 40332 1492 40352
rect 1492 40332 1544 40352
rect 1544 40332 1546 40352
rect 1490 40296 1546 40332
rect 1398 39616 1454 39672
rect 1398 39072 1454 39128
rect 1398 38528 1454 38584
rect 1398 37984 1454 38040
rect 1398 37440 1454 37496
rect 1398 36896 1454 36952
rect 1398 36352 1454 36408
rect 1398 35808 1454 35864
rect 1398 35264 1454 35320
rect 1398 34720 1454 34776
rect 1398 34176 1454 34232
rect 1398 33632 1454 33688
rect 1398 32952 1454 33008
rect 1398 32408 1454 32464
rect 1306 31864 1362 31920
rect 1398 31320 1454 31376
rect 1306 30776 1362 30832
rect 2778 62736 2834 62792
rect 2588 62586 2644 62588
rect 2668 62586 2724 62588
rect 2748 62586 2804 62588
rect 2828 62586 2884 62588
rect 2588 62534 2634 62586
rect 2634 62534 2644 62586
rect 2668 62534 2698 62586
rect 2698 62534 2710 62586
rect 2710 62534 2724 62586
rect 2748 62534 2762 62586
rect 2762 62534 2774 62586
rect 2774 62534 2804 62586
rect 2828 62534 2838 62586
rect 2838 62534 2884 62586
rect 2588 62532 2644 62534
rect 2668 62532 2724 62534
rect 2748 62532 2804 62534
rect 2828 62532 2884 62534
rect 4219 74010 4275 74012
rect 4299 74010 4355 74012
rect 4379 74010 4435 74012
rect 4459 74010 4515 74012
rect 4219 73958 4265 74010
rect 4265 73958 4275 74010
rect 4299 73958 4329 74010
rect 4329 73958 4341 74010
rect 4341 73958 4355 74010
rect 4379 73958 4393 74010
rect 4393 73958 4405 74010
rect 4405 73958 4435 74010
rect 4459 73958 4469 74010
rect 4469 73958 4515 74010
rect 4219 73956 4275 73958
rect 4299 73956 4355 73958
rect 4379 73956 4435 73958
rect 4459 73956 4515 73958
rect 4219 72922 4275 72924
rect 4299 72922 4355 72924
rect 4379 72922 4435 72924
rect 4459 72922 4515 72924
rect 4219 72870 4265 72922
rect 4265 72870 4275 72922
rect 4299 72870 4329 72922
rect 4329 72870 4341 72922
rect 4341 72870 4355 72922
rect 4379 72870 4393 72922
rect 4393 72870 4405 72922
rect 4405 72870 4435 72922
rect 4459 72870 4469 72922
rect 4469 72870 4515 72922
rect 4219 72868 4275 72870
rect 4299 72868 4355 72870
rect 4379 72868 4435 72870
rect 4459 72868 4515 72870
rect 4219 71834 4275 71836
rect 4299 71834 4355 71836
rect 4379 71834 4435 71836
rect 4459 71834 4515 71836
rect 4219 71782 4265 71834
rect 4265 71782 4275 71834
rect 4299 71782 4329 71834
rect 4329 71782 4341 71834
rect 4341 71782 4355 71834
rect 4379 71782 4393 71834
rect 4393 71782 4405 71834
rect 4405 71782 4435 71834
rect 4459 71782 4469 71834
rect 4469 71782 4515 71834
rect 4219 71780 4275 71782
rect 4299 71780 4355 71782
rect 4379 71780 4435 71782
rect 4459 71780 4515 71782
rect 3882 66544 3938 66600
rect 4219 70746 4275 70748
rect 4299 70746 4355 70748
rect 4379 70746 4435 70748
rect 4459 70746 4515 70748
rect 4219 70694 4265 70746
rect 4265 70694 4275 70746
rect 4299 70694 4329 70746
rect 4329 70694 4341 70746
rect 4341 70694 4355 70746
rect 4379 70694 4393 70746
rect 4393 70694 4405 70746
rect 4405 70694 4435 70746
rect 4459 70694 4469 70746
rect 4469 70694 4515 70746
rect 4219 70692 4275 70694
rect 4299 70692 4355 70694
rect 4379 70692 4435 70694
rect 4459 70692 4515 70694
rect 4219 69658 4275 69660
rect 4299 69658 4355 69660
rect 4379 69658 4435 69660
rect 4459 69658 4515 69660
rect 4219 69606 4265 69658
rect 4265 69606 4275 69658
rect 4299 69606 4329 69658
rect 4329 69606 4341 69658
rect 4341 69606 4355 69658
rect 4379 69606 4393 69658
rect 4393 69606 4405 69658
rect 4405 69606 4435 69658
rect 4459 69606 4469 69658
rect 4469 69606 4515 69658
rect 4219 69604 4275 69606
rect 4299 69604 4355 69606
rect 4379 69604 4435 69606
rect 4459 69604 4515 69606
rect 4219 68570 4275 68572
rect 4299 68570 4355 68572
rect 4379 68570 4435 68572
rect 4459 68570 4515 68572
rect 4219 68518 4265 68570
rect 4265 68518 4275 68570
rect 4299 68518 4329 68570
rect 4329 68518 4341 68570
rect 4341 68518 4355 68570
rect 4379 68518 4393 68570
rect 4393 68518 4405 68570
rect 4405 68518 4435 68570
rect 4459 68518 4469 68570
rect 4469 68518 4515 68570
rect 4219 68516 4275 68518
rect 4299 68516 4355 68518
rect 4379 68516 4435 68518
rect 4459 68516 4515 68518
rect 4219 67482 4275 67484
rect 4299 67482 4355 67484
rect 4379 67482 4435 67484
rect 4459 67482 4515 67484
rect 4219 67430 4265 67482
rect 4265 67430 4275 67482
rect 4299 67430 4329 67482
rect 4329 67430 4341 67482
rect 4341 67430 4355 67482
rect 4379 67430 4393 67482
rect 4393 67430 4405 67482
rect 4405 67430 4435 67482
rect 4459 67430 4469 67482
rect 4469 67430 4515 67482
rect 4219 67428 4275 67430
rect 4299 67428 4355 67430
rect 4379 67428 4435 67430
rect 4459 67428 4515 67430
rect 3882 66272 3938 66328
rect 2588 61498 2644 61500
rect 2668 61498 2724 61500
rect 2748 61498 2804 61500
rect 2828 61498 2884 61500
rect 2588 61446 2634 61498
rect 2634 61446 2644 61498
rect 2668 61446 2698 61498
rect 2698 61446 2710 61498
rect 2710 61446 2724 61498
rect 2748 61446 2762 61498
rect 2762 61446 2774 61498
rect 2774 61446 2804 61498
rect 2828 61446 2838 61498
rect 2838 61446 2884 61498
rect 2588 61444 2644 61446
rect 2668 61444 2724 61446
rect 2748 61444 2804 61446
rect 2828 61444 2884 61446
rect 2588 60410 2644 60412
rect 2668 60410 2724 60412
rect 2748 60410 2804 60412
rect 2828 60410 2884 60412
rect 2588 60358 2634 60410
rect 2634 60358 2644 60410
rect 2668 60358 2698 60410
rect 2698 60358 2710 60410
rect 2710 60358 2724 60410
rect 2748 60358 2762 60410
rect 2762 60358 2774 60410
rect 2774 60358 2804 60410
rect 2828 60358 2838 60410
rect 2838 60358 2884 60410
rect 2588 60356 2644 60358
rect 2668 60356 2724 60358
rect 2748 60356 2804 60358
rect 2828 60356 2884 60358
rect 2588 59322 2644 59324
rect 2668 59322 2724 59324
rect 2748 59322 2804 59324
rect 2828 59322 2884 59324
rect 2588 59270 2634 59322
rect 2634 59270 2644 59322
rect 2668 59270 2698 59322
rect 2698 59270 2710 59322
rect 2710 59270 2724 59322
rect 2748 59270 2762 59322
rect 2762 59270 2774 59322
rect 2774 59270 2804 59322
rect 2828 59270 2838 59322
rect 2838 59270 2884 59322
rect 2588 59268 2644 59270
rect 2668 59268 2724 59270
rect 2748 59268 2804 59270
rect 2828 59268 2884 59270
rect 2588 58234 2644 58236
rect 2668 58234 2724 58236
rect 2748 58234 2804 58236
rect 2828 58234 2884 58236
rect 2588 58182 2634 58234
rect 2634 58182 2644 58234
rect 2668 58182 2698 58234
rect 2698 58182 2710 58234
rect 2710 58182 2724 58234
rect 2748 58182 2762 58234
rect 2762 58182 2774 58234
rect 2774 58182 2804 58234
rect 2828 58182 2838 58234
rect 2838 58182 2884 58234
rect 2588 58180 2644 58182
rect 2668 58180 2724 58182
rect 2748 58180 2804 58182
rect 2828 58180 2884 58182
rect 2778 57432 2834 57488
rect 2588 57146 2644 57148
rect 2668 57146 2724 57148
rect 2748 57146 2804 57148
rect 2828 57146 2884 57148
rect 2588 57094 2634 57146
rect 2634 57094 2644 57146
rect 2668 57094 2698 57146
rect 2698 57094 2710 57146
rect 2710 57094 2724 57146
rect 2748 57094 2762 57146
rect 2762 57094 2774 57146
rect 2774 57094 2804 57146
rect 2828 57094 2838 57146
rect 2838 57094 2884 57146
rect 2588 57092 2644 57094
rect 2668 57092 2724 57094
rect 2748 57092 2804 57094
rect 2828 57092 2884 57094
rect 2588 56058 2644 56060
rect 2668 56058 2724 56060
rect 2748 56058 2804 56060
rect 2828 56058 2884 56060
rect 2588 56006 2634 56058
rect 2634 56006 2644 56058
rect 2668 56006 2698 56058
rect 2698 56006 2710 56058
rect 2710 56006 2724 56058
rect 2748 56006 2762 56058
rect 2762 56006 2774 56058
rect 2774 56006 2804 56058
rect 2828 56006 2838 56058
rect 2838 56006 2884 56058
rect 2588 56004 2644 56006
rect 2668 56004 2724 56006
rect 2748 56004 2804 56006
rect 2828 56004 2884 56006
rect 3054 56228 3110 56264
rect 3054 56208 3056 56228
rect 3056 56208 3108 56228
rect 3108 56208 3110 56228
rect 2962 55800 3018 55856
rect 2588 54970 2644 54972
rect 2668 54970 2724 54972
rect 2748 54970 2804 54972
rect 2828 54970 2884 54972
rect 2588 54918 2634 54970
rect 2634 54918 2644 54970
rect 2668 54918 2698 54970
rect 2698 54918 2710 54970
rect 2710 54918 2724 54970
rect 2748 54918 2762 54970
rect 2762 54918 2774 54970
rect 2774 54918 2804 54970
rect 2828 54918 2838 54970
rect 2838 54918 2884 54970
rect 2588 54916 2644 54918
rect 2668 54916 2724 54918
rect 2748 54916 2804 54918
rect 2828 54916 2884 54918
rect 2962 54712 3018 54768
rect 2588 53882 2644 53884
rect 2668 53882 2724 53884
rect 2748 53882 2804 53884
rect 2828 53882 2884 53884
rect 2588 53830 2634 53882
rect 2634 53830 2644 53882
rect 2668 53830 2698 53882
rect 2698 53830 2710 53882
rect 2710 53830 2724 53882
rect 2748 53830 2762 53882
rect 2762 53830 2774 53882
rect 2774 53830 2804 53882
rect 2828 53830 2838 53882
rect 2838 53830 2884 53882
rect 2588 53828 2644 53830
rect 2668 53828 2724 53830
rect 2748 53828 2804 53830
rect 2828 53828 2884 53830
rect 2778 52944 2834 53000
rect 2588 52794 2644 52796
rect 2668 52794 2724 52796
rect 2748 52794 2804 52796
rect 2828 52794 2884 52796
rect 2588 52742 2634 52794
rect 2634 52742 2644 52794
rect 2668 52742 2698 52794
rect 2698 52742 2710 52794
rect 2710 52742 2724 52794
rect 2748 52742 2762 52794
rect 2762 52742 2774 52794
rect 2774 52742 2804 52794
rect 2828 52742 2838 52794
rect 2838 52742 2884 52794
rect 2588 52740 2644 52742
rect 2668 52740 2724 52742
rect 2748 52740 2804 52742
rect 2828 52740 2884 52742
rect 2502 52128 2558 52184
rect 2318 51584 2374 51640
rect 2410 51448 2466 51504
rect 2226 51040 2282 51096
rect 1398 30232 1454 30288
rect 1306 29688 1362 29744
rect 1398 29144 1454 29200
rect 1306 28600 1362 28656
rect 1398 28056 1454 28112
rect 1306 27512 1362 27568
rect 1950 41112 2006 41168
rect 2134 41656 2190 41712
rect 2318 41248 2374 41304
rect 2318 41112 2374 41168
rect 2778 51876 2834 51912
rect 2778 51856 2780 51876
rect 2780 51856 2832 51876
rect 2832 51856 2834 51876
rect 2588 51706 2644 51708
rect 2668 51706 2724 51708
rect 2748 51706 2804 51708
rect 2828 51706 2884 51708
rect 2588 51654 2634 51706
rect 2634 51654 2644 51706
rect 2668 51654 2698 51706
rect 2698 51654 2710 51706
rect 2710 51654 2724 51706
rect 2748 51654 2762 51706
rect 2762 51654 2774 51706
rect 2774 51654 2804 51706
rect 2828 51654 2838 51706
rect 2838 51654 2884 51706
rect 2588 51652 2644 51654
rect 2668 51652 2724 51654
rect 2748 51652 2804 51654
rect 2828 51652 2884 51654
rect 3238 53080 3294 53136
rect 2594 51312 2650 51368
rect 3146 52808 3202 52864
rect 2778 50788 2834 50824
rect 2778 50768 2780 50788
rect 2780 50768 2832 50788
rect 2832 50768 2834 50788
rect 2588 50618 2644 50620
rect 2668 50618 2724 50620
rect 2748 50618 2804 50620
rect 2828 50618 2884 50620
rect 2588 50566 2634 50618
rect 2634 50566 2644 50618
rect 2668 50566 2698 50618
rect 2698 50566 2710 50618
rect 2710 50566 2724 50618
rect 2748 50566 2762 50618
rect 2762 50566 2774 50618
rect 2774 50566 2804 50618
rect 2828 50566 2838 50618
rect 2838 50566 2884 50618
rect 2588 50564 2644 50566
rect 2668 50564 2724 50566
rect 2748 50564 2804 50566
rect 2828 50564 2884 50566
rect 2502 50224 2558 50280
rect 2588 49530 2644 49532
rect 2668 49530 2724 49532
rect 2748 49530 2804 49532
rect 2828 49530 2884 49532
rect 2588 49478 2634 49530
rect 2634 49478 2644 49530
rect 2668 49478 2698 49530
rect 2698 49478 2710 49530
rect 2710 49478 2724 49530
rect 2748 49478 2762 49530
rect 2762 49478 2774 49530
rect 2774 49478 2804 49530
rect 2828 49478 2838 49530
rect 2838 49478 2884 49530
rect 2588 49476 2644 49478
rect 2668 49476 2724 49478
rect 2748 49476 2804 49478
rect 2828 49476 2884 49478
rect 2588 48442 2644 48444
rect 2668 48442 2724 48444
rect 2748 48442 2804 48444
rect 2828 48442 2884 48444
rect 2588 48390 2634 48442
rect 2634 48390 2644 48442
rect 2668 48390 2698 48442
rect 2698 48390 2710 48442
rect 2710 48390 2724 48442
rect 2748 48390 2762 48442
rect 2762 48390 2774 48442
rect 2774 48390 2804 48442
rect 2828 48390 2838 48442
rect 2838 48390 2884 48442
rect 2588 48388 2644 48390
rect 2668 48388 2724 48390
rect 2748 48388 2804 48390
rect 2828 48388 2884 48390
rect 2588 47354 2644 47356
rect 2668 47354 2724 47356
rect 2748 47354 2804 47356
rect 2828 47354 2884 47356
rect 2588 47302 2634 47354
rect 2634 47302 2644 47354
rect 2668 47302 2698 47354
rect 2698 47302 2710 47354
rect 2710 47302 2724 47354
rect 2748 47302 2762 47354
rect 2762 47302 2774 47354
rect 2774 47302 2804 47354
rect 2828 47302 2838 47354
rect 2838 47302 2884 47354
rect 2588 47300 2644 47302
rect 2668 47300 2724 47302
rect 2748 47300 2804 47302
rect 2828 47300 2884 47302
rect 2588 46266 2644 46268
rect 2668 46266 2724 46268
rect 2748 46266 2804 46268
rect 2828 46266 2884 46268
rect 2588 46214 2634 46266
rect 2634 46214 2644 46266
rect 2668 46214 2698 46266
rect 2698 46214 2710 46266
rect 2710 46214 2724 46266
rect 2748 46214 2762 46266
rect 2762 46214 2774 46266
rect 2774 46214 2804 46266
rect 2828 46214 2838 46266
rect 2838 46214 2884 46266
rect 2588 46212 2644 46214
rect 2668 46212 2724 46214
rect 2748 46212 2804 46214
rect 2828 46212 2884 46214
rect 2686 46008 2742 46064
rect 2588 45178 2644 45180
rect 2668 45178 2724 45180
rect 2748 45178 2804 45180
rect 2828 45178 2884 45180
rect 2588 45126 2634 45178
rect 2634 45126 2644 45178
rect 2668 45126 2698 45178
rect 2698 45126 2710 45178
rect 2710 45126 2724 45178
rect 2748 45126 2762 45178
rect 2762 45126 2774 45178
rect 2774 45126 2804 45178
rect 2828 45126 2838 45178
rect 2838 45126 2884 45178
rect 2588 45124 2644 45126
rect 2668 45124 2724 45126
rect 2748 45124 2804 45126
rect 2828 45124 2884 45126
rect 3238 52128 3294 52184
rect 3974 63008 4030 63064
rect 3514 52264 3570 52320
rect 3514 50768 3570 50824
rect 2588 44090 2644 44092
rect 2668 44090 2724 44092
rect 2748 44090 2804 44092
rect 2828 44090 2884 44092
rect 2588 44038 2634 44090
rect 2634 44038 2644 44090
rect 2668 44038 2698 44090
rect 2698 44038 2710 44090
rect 2710 44038 2724 44090
rect 2748 44038 2762 44090
rect 2762 44038 2774 44090
rect 2774 44038 2804 44090
rect 2828 44038 2838 44090
rect 2838 44038 2884 44090
rect 2588 44036 2644 44038
rect 2668 44036 2724 44038
rect 2748 44036 2804 44038
rect 2828 44036 2884 44038
rect 2588 43002 2644 43004
rect 2668 43002 2724 43004
rect 2748 43002 2804 43004
rect 2828 43002 2884 43004
rect 2588 42950 2634 43002
rect 2634 42950 2644 43002
rect 2668 42950 2698 43002
rect 2698 42950 2710 43002
rect 2710 42950 2724 43002
rect 2748 42950 2762 43002
rect 2762 42950 2774 43002
rect 2774 42950 2804 43002
rect 2828 42950 2838 43002
rect 2838 42950 2884 43002
rect 2588 42948 2644 42950
rect 2668 42948 2724 42950
rect 2748 42948 2804 42950
rect 2828 42948 2884 42950
rect 2588 41914 2644 41916
rect 2668 41914 2724 41916
rect 2748 41914 2804 41916
rect 2828 41914 2884 41916
rect 2588 41862 2634 41914
rect 2634 41862 2644 41914
rect 2668 41862 2698 41914
rect 2698 41862 2710 41914
rect 2710 41862 2724 41914
rect 2748 41862 2762 41914
rect 2762 41862 2774 41914
rect 2774 41862 2804 41914
rect 2828 41862 2838 41914
rect 2838 41862 2884 41914
rect 2588 41860 2644 41862
rect 2668 41860 2724 41862
rect 2748 41860 2804 41862
rect 2828 41860 2884 41862
rect 2502 41520 2558 41576
rect 2502 41112 2558 41168
rect 2778 41112 2834 41168
rect 2588 40826 2644 40828
rect 2668 40826 2724 40828
rect 2748 40826 2804 40828
rect 2828 40826 2884 40828
rect 2588 40774 2634 40826
rect 2634 40774 2644 40826
rect 2668 40774 2698 40826
rect 2698 40774 2710 40826
rect 2710 40774 2724 40826
rect 2748 40774 2762 40826
rect 2762 40774 2774 40826
rect 2774 40774 2804 40826
rect 2828 40774 2838 40826
rect 2838 40774 2884 40826
rect 2588 40772 2644 40774
rect 2668 40772 2724 40774
rect 2748 40772 2804 40774
rect 2828 40772 2884 40774
rect 2594 40044 2650 40080
rect 2594 40024 2596 40044
rect 2596 40024 2648 40044
rect 2648 40024 2650 40044
rect 2588 39738 2644 39740
rect 2668 39738 2724 39740
rect 2748 39738 2804 39740
rect 2828 39738 2884 39740
rect 2588 39686 2634 39738
rect 2634 39686 2644 39738
rect 2668 39686 2698 39738
rect 2698 39686 2710 39738
rect 2710 39686 2724 39738
rect 2748 39686 2762 39738
rect 2762 39686 2774 39738
rect 2774 39686 2804 39738
rect 2828 39686 2838 39738
rect 2838 39686 2884 39738
rect 2588 39684 2644 39686
rect 2668 39684 2724 39686
rect 2748 39684 2804 39686
rect 2828 39684 2884 39686
rect 2588 38650 2644 38652
rect 2668 38650 2724 38652
rect 2748 38650 2804 38652
rect 2828 38650 2884 38652
rect 2588 38598 2634 38650
rect 2634 38598 2644 38650
rect 2668 38598 2698 38650
rect 2698 38598 2710 38650
rect 2710 38598 2724 38650
rect 2748 38598 2762 38650
rect 2762 38598 2774 38650
rect 2774 38598 2804 38650
rect 2828 38598 2838 38650
rect 2838 38598 2884 38650
rect 2588 38596 2644 38598
rect 2668 38596 2724 38598
rect 2748 38596 2804 38598
rect 2828 38596 2884 38598
rect 2588 37562 2644 37564
rect 2668 37562 2724 37564
rect 2748 37562 2804 37564
rect 2828 37562 2884 37564
rect 2588 37510 2634 37562
rect 2634 37510 2644 37562
rect 2668 37510 2698 37562
rect 2698 37510 2710 37562
rect 2710 37510 2724 37562
rect 2748 37510 2762 37562
rect 2762 37510 2774 37562
rect 2774 37510 2804 37562
rect 2828 37510 2838 37562
rect 2838 37510 2884 37562
rect 2588 37508 2644 37510
rect 2668 37508 2724 37510
rect 2748 37508 2804 37510
rect 2828 37508 2884 37510
rect 2588 36474 2644 36476
rect 2668 36474 2724 36476
rect 2748 36474 2804 36476
rect 2828 36474 2884 36476
rect 2588 36422 2634 36474
rect 2634 36422 2644 36474
rect 2668 36422 2698 36474
rect 2698 36422 2710 36474
rect 2710 36422 2724 36474
rect 2748 36422 2762 36474
rect 2762 36422 2774 36474
rect 2774 36422 2804 36474
rect 2828 36422 2838 36474
rect 2838 36422 2884 36474
rect 2588 36420 2644 36422
rect 2668 36420 2724 36422
rect 2748 36420 2804 36422
rect 2828 36420 2884 36422
rect 2588 35386 2644 35388
rect 2668 35386 2724 35388
rect 2748 35386 2804 35388
rect 2828 35386 2884 35388
rect 2588 35334 2634 35386
rect 2634 35334 2644 35386
rect 2668 35334 2698 35386
rect 2698 35334 2710 35386
rect 2710 35334 2724 35386
rect 2748 35334 2762 35386
rect 2762 35334 2774 35386
rect 2774 35334 2804 35386
rect 2828 35334 2838 35386
rect 2838 35334 2884 35386
rect 2588 35332 2644 35334
rect 2668 35332 2724 35334
rect 2748 35332 2804 35334
rect 2828 35332 2884 35334
rect 2588 34298 2644 34300
rect 2668 34298 2724 34300
rect 2748 34298 2804 34300
rect 2828 34298 2884 34300
rect 2588 34246 2634 34298
rect 2634 34246 2644 34298
rect 2668 34246 2698 34298
rect 2698 34246 2710 34298
rect 2710 34246 2724 34298
rect 2748 34246 2762 34298
rect 2762 34246 2774 34298
rect 2774 34246 2804 34298
rect 2828 34246 2838 34298
rect 2838 34246 2884 34298
rect 2588 34244 2644 34246
rect 2668 34244 2724 34246
rect 2748 34244 2804 34246
rect 2828 34244 2884 34246
rect 2588 33210 2644 33212
rect 2668 33210 2724 33212
rect 2748 33210 2804 33212
rect 2828 33210 2884 33212
rect 2588 33158 2634 33210
rect 2634 33158 2644 33210
rect 2668 33158 2698 33210
rect 2698 33158 2710 33210
rect 2710 33158 2724 33210
rect 2748 33158 2762 33210
rect 2762 33158 2774 33210
rect 2774 33158 2804 33210
rect 2828 33158 2838 33210
rect 2838 33158 2884 33210
rect 2588 33156 2644 33158
rect 2668 33156 2724 33158
rect 2748 33156 2804 33158
rect 2828 33156 2884 33158
rect 2588 32122 2644 32124
rect 2668 32122 2724 32124
rect 2748 32122 2804 32124
rect 2828 32122 2884 32124
rect 2588 32070 2634 32122
rect 2634 32070 2644 32122
rect 2668 32070 2698 32122
rect 2698 32070 2710 32122
rect 2710 32070 2724 32122
rect 2748 32070 2762 32122
rect 2762 32070 2774 32122
rect 2774 32070 2804 32122
rect 2828 32070 2838 32122
rect 2838 32070 2884 32122
rect 2588 32068 2644 32070
rect 2668 32068 2724 32070
rect 2748 32068 2804 32070
rect 2828 32068 2884 32070
rect 2588 31034 2644 31036
rect 2668 31034 2724 31036
rect 2748 31034 2804 31036
rect 2828 31034 2884 31036
rect 2588 30982 2634 31034
rect 2634 30982 2644 31034
rect 2668 30982 2698 31034
rect 2698 30982 2710 31034
rect 2710 30982 2724 31034
rect 2748 30982 2762 31034
rect 2762 30982 2774 31034
rect 2774 30982 2804 31034
rect 2828 30982 2838 31034
rect 2838 30982 2884 31034
rect 2588 30980 2644 30982
rect 2668 30980 2724 30982
rect 2748 30980 2804 30982
rect 2828 30980 2884 30982
rect 3238 45464 3294 45520
rect 3238 45056 3294 45112
rect 3054 40024 3110 40080
rect 2588 29946 2644 29948
rect 2668 29946 2724 29948
rect 2748 29946 2804 29948
rect 2828 29946 2884 29948
rect 2588 29894 2634 29946
rect 2634 29894 2644 29946
rect 2668 29894 2698 29946
rect 2698 29894 2710 29946
rect 2710 29894 2724 29946
rect 2748 29894 2762 29946
rect 2762 29894 2774 29946
rect 2774 29894 2804 29946
rect 2828 29894 2838 29946
rect 2838 29894 2884 29946
rect 2588 29892 2644 29894
rect 2668 29892 2724 29894
rect 2748 29892 2804 29894
rect 2828 29892 2884 29894
rect 2588 28858 2644 28860
rect 2668 28858 2724 28860
rect 2748 28858 2804 28860
rect 2828 28858 2884 28860
rect 2588 28806 2634 28858
rect 2634 28806 2644 28858
rect 2668 28806 2698 28858
rect 2698 28806 2710 28858
rect 2710 28806 2724 28858
rect 2748 28806 2762 28858
rect 2762 28806 2774 28858
rect 2774 28806 2804 28858
rect 2828 28806 2838 28858
rect 2838 28806 2884 28858
rect 2588 28804 2644 28806
rect 2668 28804 2724 28806
rect 2748 28804 2804 28806
rect 2828 28804 2884 28806
rect 2588 27770 2644 27772
rect 2668 27770 2724 27772
rect 2748 27770 2804 27772
rect 2828 27770 2884 27772
rect 2588 27718 2634 27770
rect 2634 27718 2644 27770
rect 2668 27718 2698 27770
rect 2698 27718 2710 27770
rect 2710 27718 2724 27770
rect 2748 27718 2762 27770
rect 2762 27718 2774 27770
rect 2774 27718 2804 27770
rect 2828 27718 2838 27770
rect 2838 27718 2884 27770
rect 2588 27716 2644 27718
rect 2668 27716 2724 27718
rect 2748 27716 2804 27718
rect 2828 27716 2884 27718
rect 1950 26968 2006 27024
rect 1950 26308 2006 26344
rect 1950 26288 1952 26308
rect 1952 26288 2004 26308
rect 2004 26288 2006 26308
rect 1950 25744 2006 25800
rect 1950 25220 2006 25256
rect 1950 25200 1952 25220
rect 1952 25200 2004 25220
rect 2004 25200 2006 25220
rect 1950 24656 2006 24712
rect 1950 24132 2006 24168
rect 1950 24112 1952 24132
rect 1952 24112 2004 24132
rect 2004 24112 2006 24132
rect 1490 21412 1546 21448
rect 1490 21392 1492 21412
rect 1492 21392 1544 21412
rect 1544 21392 1546 21412
rect 1490 20848 1546 20904
rect 1490 20324 1546 20360
rect 1490 20304 1492 20324
rect 1492 20304 1544 20324
rect 1544 20304 1546 20324
rect 1490 19660 1492 19680
rect 1492 19660 1544 19680
rect 1544 19660 1546 19680
rect 1490 19624 1546 19660
rect 1490 19116 1492 19136
rect 1492 19116 1544 19136
rect 1544 19116 1546 19136
rect 1490 19080 1546 19116
rect 1858 23568 1914 23624
rect 1950 23044 2006 23080
rect 1950 23024 1952 23044
rect 1952 23024 2004 23044
rect 2004 23024 2006 23044
rect 1950 22480 2006 22536
rect 1950 21972 1952 21992
rect 1952 21972 2004 21992
rect 2004 21972 2006 21992
rect 1950 21936 2006 21972
rect 1490 18572 1492 18592
rect 1492 18572 1544 18592
rect 1544 18572 1546 18592
rect 1490 18536 1546 18572
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 1490 17484 1492 17504
rect 1492 17484 1544 17504
rect 1544 17484 1546 17504
rect 1490 17448 1546 17484
rect 1490 16940 1492 16960
rect 1492 16940 1544 16960
rect 1544 16940 1546 16960
rect 1490 16904 1546 16940
rect 1490 16396 1492 16416
rect 1492 16396 1544 16416
rect 1544 16396 1546 16416
rect 1490 16360 1546 16396
rect 1490 15852 1492 15872
rect 1492 15852 1544 15872
rect 1544 15852 1546 15872
rect 1490 15816 1546 15852
rect 1490 15308 1492 15328
rect 1492 15308 1544 15328
rect 1544 15308 1546 15328
rect 1490 15272 1546 15308
rect 1490 14764 1492 14784
rect 1492 14764 1544 14784
rect 1544 14764 1546 14784
rect 1490 14728 1546 14764
rect 1490 14220 1492 14240
rect 1492 14220 1544 14240
rect 1544 14220 1546 14240
rect 1490 14184 1546 14220
rect 1490 13676 1492 13696
rect 1492 13676 1544 13696
rect 1544 13676 1546 13696
rect 1490 13640 1546 13676
rect 1490 12960 1546 13016
rect 1490 12416 1546 12472
rect 1490 11872 1546 11928
rect 1490 11328 1546 11384
rect 1490 10784 1546 10840
rect 1490 10240 1546 10296
rect 1490 9696 1546 9752
rect 1490 8608 1546 8664
rect 1398 8064 1454 8120
rect 1490 7520 1546 7576
rect 1306 6296 1362 6352
rect 1490 5752 1546 5808
rect 2588 26682 2644 26684
rect 2668 26682 2724 26684
rect 2748 26682 2804 26684
rect 2828 26682 2884 26684
rect 2588 26630 2634 26682
rect 2634 26630 2644 26682
rect 2668 26630 2698 26682
rect 2698 26630 2710 26682
rect 2710 26630 2724 26682
rect 2748 26630 2762 26682
rect 2762 26630 2774 26682
rect 2774 26630 2804 26682
rect 2828 26630 2838 26682
rect 2838 26630 2884 26682
rect 2588 26628 2644 26630
rect 2668 26628 2724 26630
rect 2748 26628 2804 26630
rect 2828 26628 2884 26630
rect 2588 25594 2644 25596
rect 2668 25594 2724 25596
rect 2748 25594 2804 25596
rect 2828 25594 2884 25596
rect 2588 25542 2634 25594
rect 2634 25542 2644 25594
rect 2668 25542 2698 25594
rect 2698 25542 2710 25594
rect 2710 25542 2724 25594
rect 2748 25542 2762 25594
rect 2762 25542 2774 25594
rect 2774 25542 2804 25594
rect 2828 25542 2838 25594
rect 2838 25542 2884 25594
rect 2588 25540 2644 25542
rect 2668 25540 2724 25542
rect 2748 25540 2804 25542
rect 2828 25540 2884 25542
rect 2588 24506 2644 24508
rect 2668 24506 2724 24508
rect 2748 24506 2804 24508
rect 2828 24506 2884 24508
rect 2588 24454 2634 24506
rect 2634 24454 2644 24506
rect 2668 24454 2698 24506
rect 2698 24454 2710 24506
rect 2710 24454 2724 24506
rect 2748 24454 2762 24506
rect 2762 24454 2774 24506
rect 2774 24454 2804 24506
rect 2828 24454 2838 24506
rect 2838 24454 2884 24506
rect 2588 24452 2644 24454
rect 2668 24452 2724 24454
rect 2748 24452 2804 24454
rect 2828 24452 2884 24454
rect 3698 48592 3754 48648
rect 3698 48320 3754 48376
rect 3606 46280 3662 46336
rect 4219 66394 4275 66396
rect 4299 66394 4355 66396
rect 4379 66394 4435 66396
rect 4459 66394 4515 66396
rect 4219 66342 4265 66394
rect 4265 66342 4275 66394
rect 4299 66342 4329 66394
rect 4329 66342 4341 66394
rect 4341 66342 4355 66394
rect 4379 66342 4393 66394
rect 4393 66342 4405 66394
rect 4405 66342 4435 66394
rect 4459 66342 4469 66394
rect 4469 66342 4515 66394
rect 4219 66340 4275 66342
rect 4299 66340 4355 66342
rect 4379 66340 4435 66342
rect 4459 66340 4515 66342
rect 4219 65306 4275 65308
rect 4299 65306 4355 65308
rect 4379 65306 4435 65308
rect 4459 65306 4515 65308
rect 4219 65254 4265 65306
rect 4265 65254 4275 65306
rect 4299 65254 4329 65306
rect 4329 65254 4341 65306
rect 4341 65254 4355 65306
rect 4379 65254 4393 65306
rect 4393 65254 4405 65306
rect 4405 65254 4435 65306
rect 4459 65254 4469 65306
rect 4469 65254 4515 65306
rect 4219 65252 4275 65254
rect 4299 65252 4355 65254
rect 4379 65252 4435 65254
rect 4459 65252 4515 65254
rect 4219 64218 4275 64220
rect 4299 64218 4355 64220
rect 4379 64218 4435 64220
rect 4459 64218 4515 64220
rect 4219 64166 4265 64218
rect 4265 64166 4275 64218
rect 4299 64166 4329 64218
rect 4329 64166 4341 64218
rect 4341 64166 4355 64218
rect 4379 64166 4393 64218
rect 4393 64166 4405 64218
rect 4405 64166 4435 64218
rect 4459 64166 4469 64218
rect 4469 64166 4515 64218
rect 4219 64164 4275 64166
rect 4299 64164 4355 64166
rect 4379 64164 4435 64166
rect 4459 64164 4515 64166
rect 4219 63130 4275 63132
rect 4299 63130 4355 63132
rect 4379 63130 4435 63132
rect 4459 63130 4515 63132
rect 4219 63078 4265 63130
rect 4265 63078 4275 63130
rect 4299 63078 4329 63130
rect 4329 63078 4341 63130
rect 4341 63078 4355 63130
rect 4379 63078 4393 63130
rect 4393 63078 4405 63130
rect 4405 63078 4435 63130
rect 4459 63078 4469 63130
rect 4469 63078 4515 63130
rect 4219 63076 4275 63078
rect 4299 63076 4355 63078
rect 4379 63076 4435 63078
rect 4459 63076 4515 63078
rect 4219 62042 4275 62044
rect 4299 62042 4355 62044
rect 4379 62042 4435 62044
rect 4459 62042 4515 62044
rect 4219 61990 4265 62042
rect 4265 61990 4275 62042
rect 4299 61990 4329 62042
rect 4329 61990 4341 62042
rect 4341 61990 4355 62042
rect 4379 61990 4393 62042
rect 4393 61990 4405 62042
rect 4405 61990 4435 62042
rect 4459 61990 4469 62042
rect 4469 61990 4515 62042
rect 4219 61988 4275 61990
rect 4299 61988 4355 61990
rect 4379 61988 4435 61990
rect 4459 61988 4515 61990
rect 4219 60954 4275 60956
rect 4299 60954 4355 60956
rect 4379 60954 4435 60956
rect 4459 60954 4515 60956
rect 4219 60902 4265 60954
rect 4265 60902 4275 60954
rect 4299 60902 4329 60954
rect 4329 60902 4341 60954
rect 4341 60902 4355 60954
rect 4379 60902 4393 60954
rect 4393 60902 4405 60954
rect 4405 60902 4435 60954
rect 4459 60902 4469 60954
rect 4469 60902 4515 60954
rect 4219 60900 4275 60902
rect 4299 60900 4355 60902
rect 4379 60900 4435 60902
rect 4459 60900 4515 60902
rect 4219 59866 4275 59868
rect 4299 59866 4355 59868
rect 4379 59866 4435 59868
rect 4459 59866 4515 59868
rect 4219 59814 4265 59866
rect 4265 59814 4275 59866
rect 4299 59814 4329 59866
rect 4329 59814 4341 59866
rect 4341 59814 4355 59866
rect 4379 59814 4393 59866
rect 4393 59814 4405 59866
rect 4405 59814 4435 59866
rect 4459 59814 4469 59866
rect 4469 59814 4515 59866
rect 4219 59812 4275 59814
rect 4299 59812 4355 59814
rect 4379 59812 4435 59814
rect 4459 59812 4515 59814
rect 4219 58778 4275 58780
rect 4299 58778 4355 58780
rect 4379 58778 4435 58780
rect 4459 58778 4515 58780
rect 4219 58726 4265 58778
rect 4265 58726 4275 58778
rect 4299 58726 4329 58778
rect 4329 58726 4341 58778
rect 4341 58726 4355 58778
rect 4379 58726 4393 58778
rect 4393 58726 4405 58778
rect 4405 58726 4435 58778
rect 4459 58726 4469 58778
rect 4469 58726 4515 58778
rect 4219 58724 4275 58726
rect 4299 58724 4355 58726
rect 4379 58724 4435 58726
rect 4459 58724 4515 58726
rect 4219 57690 4275 57692
rect 4299 57690 4355 57692
rect 4379 57690 4435 57692
rect 4459 57690 4515 57692
rect 4219 57638 4265 57690
rect 4265 57638 4275 57690
rect 4299 57638 4329 57690
rect 4329 57638 4341 57690
rect 4341 57638 4355 57690
rect 4379 57638 4393 57690
rect 4393 57638 4405 57690
rect 4405 57638 4435 57690
rect 4459 57638 4469 57690
rect 4469 57638 4515 57690
rect 4219 57636 4275 57638
rect 4299 57636 4355 57638
rect 4379 57636 4435 57638
rect 4459 57636 4515 57638
rect 4219 56602 4275 56604
rect 4299 56602 4355 56604
rect 4379 56602 4435 56604
rect 4459 56602 4515 56604
rect 4219 56550 4265 56602
rect 4265 56550 4275 56602
rect 4299 56550 4329 56602
rect 4329 56550 4341 56602
rect 4341 56550 4355 56602
rect 4379 56550 4393 56602
rect 4393 56550 4405 56602
rect 4405 56550 4435 56602
rect 4459 56550 4469 56602
rect 4469 56550 4515 56602
rect 4219 56548 4275 56550
rect 4299 56548 4355 56550
rect 4379 56548 4435 56550
rect 4459 56548 4515 56550
rect 3974 56344 4030 56400
rect 3974 55256 4030 55312
rect 4219 55514 4275 55516
rect 4299 55514 4355 55516
rect 4379 55514 4435 55516
rect 4459 55514 4515 55516
rect 4219 55462 4265 55514
rect 4265 55462 4275 55514
rect 4299 55462 4329 55514
rect 4329 55462 4341 55514
rect 4341 55462 4355 55514
rect 4379 55462 4393 55514
rect 4393 55462 4405 55514
rect 4405 55462 4435 55514
rect 4459 55462 4469 55514
rect 4469 55462 4515 55514
rect 4219 55460 4275 55462
rect 4299 55460 4355 55462
rect 4379 55460 4435 55462
rect 4459 55460 4515 55462
rect 4219 54426 4275 54428
rect 4299 54426 4355 54428
rect 4379 54426 4435 54428
rect 4459 54426 4515 54428
rect 4219 54374 4265 54426
rect 4265 54374 4275 54426
rect 4299 54374 4329 54426
rect 4329 54374 4341 54426
rect 4341 54374 4355 54426
rect 4379 54374 4393 54426
rect 4393 54374 4405 54426
rect 4405 54374 4435 54426
rect 4459 54374 4469 54426
rect 4469 54374 4515 54426
rect 4219 54372 4275 54374
rect 4299 54372 4355 54374
rect 4379 54372 4435 54374
rect 4459 54372 4515 54374
rect 4219 53338 4275 53340
rect 4299 53338 4355 53340
rect 4379 53338 4435 53340
rect 4459 53338 4515 53340
rect 4219 53286 4265 53338
rect 4265 53286 4275 53338
rect 4299 53286 4329 53338
rect 4329 53286 4341 53338
rect 4341 53286 4355 53338
rect 4379 53286 4393 53338
rect 4393 53286 4405 53338
rect 4405 53286 4435 53338
rect 4459 53286 4469 53338
rect 4469 53286 4515 53338
rect 4219 53284 4275 53286
rect 4299 53284 4355 53286
rect 4379 53284 4435 53286
rect 4459 53284 4515 53286
rect 4219 52250 4275 52252
rect 4299 52250 4355 52252
rect 4379 52250 4435 52252
rect 4459 52250 4515 52252
rect 4219 52198 4265 52250
rect 4265 52198 4275 52250
rect 4299 52198 4329 52250
rect 4329 52198 4341 52250
rect 4341 52198 4355 52250
rect 4379 52198 4393 52250
rect 4393 52198 4405 52250
rect 4405 52198 4435 52250
rect 4459 52198 4469 52250
rect 4469 52198 4515 52250
rect 4219 52196 4275 52198
rect 4299 52196 4355 52198
rect 4379 52196 4435 52198
rect 4459 52196 4515 52198
rect 3974 51032 4030 51088
rect 4219 51162 4275 51164
rect 4299 51162 4355 51164
rect 4379 51162 4435 51164
rect 4459 51162 4515 51164
rect 4219 51110 4265 51162
rect 4265 51110 4275 51162
rect 4299 51110 4329 51162
rect 4329 51110 4341 51162
rect 4341 51110 4355 51162
rect 4379 51110 4393 51162
rect 4393 51110 4405 51162
rect 4405 51110 4435 51162
rect 4459 51110 4469 51162
rect 4469 51110 4515 51162
rect 4219 51108 4275 51110
rect 4299 51108 4355 51110
rect 4379 51108 4435 51110
rect 4459 51108 4515 51110
rect 4219 50074 4275 50076
rect 4299 50074 4355 50076
rect 4379 50074 4435 50076
rect 4459 50074 4515 50076
rect 4219 50022 4265 50074
rect 4265 50022 4275 50074
rect 4299 50022 4329 50074
rect 4329 50022 4341 50074
rect 4341 50022 4355 50074
rect 4379 50022 4393 50074
rect 4393 50022 4405 50074
rect 4405 50022 4435 50074
rect 4459 50022 4469 50074
rect 4469 50022 4515 50074
rect 4219 50020 4275 50022
rect 4299 50020 4355 50022
rect 4379 50020 4435 50022
rect 4459 50020 4515 50022
rect 4219 48986 4275 48988
rect 4299 48986 4355 48988
rect 4379 48986 4435 48988
rect 4459 48986 4515 48988
rect 4219 48934 4265 48986
rect 4265 48934 4275 48986
rect 4299 48934 4329 48986
rect 4329 48934 4341 48986
rect 4341 48934 4355 48986
rect 4379 48934 4393 48986
rect 4393 48934 4405 48986
rect 4405 48934 4435 48986
rect 4459 48934 4469 48986
rect 4469 48934 4515 48986
rect 4219 48932 4275 48934
rect 4299 48932 4355 48934
rect 4379 48932 4435 48934
rect 4459 48932 4515 48934
rect 4219 47898 4275 47900
rect 4299 47898 4355 47900
rect 4379 47898 4435 47900
rect 4459 47898 4515 47900
rect 4219 47846 4265 47898
rect 4265 47846 4275 47898
rect 4299 47846 4329 47898
rect 4329 47846 4341 47898
rect 4341 47846 4355 47898
rect 4379 47846 4393 47898
rect 4393 47846 4405 47898
rect 4405 47846 4435 47898
rect 4459 47846 4469 47898
rect 4469 47846 4515 47898
rect 4219 47844 4275 47846
rect 4299 47844 4355 47846
rect 4379 47844 4435 47846
rect 4459 47844 4515 47846
rect 3974 47096 4030 47152
rect 4219 46810 4275 46812
rect 4299 46810 4355 46812
rect 4379 46810 4435 46812
rect 4459 46810 4515 46812
rect 4219 46758 4265 46810
rect 4265 46758 4275 46810
rect 4299 46758 4329 46810
rect 4329 46758 4341 46810
rect 4341 46758 4355 46810
rect 4379 46758 4393 46810
rect 4393 46758 4405 46810
rect 4405 46758 4435 46810
rect 4459 46758 4469 46810
rect 4469 46758 4515 46810
rect 4219 46756 4275 46758
rect 4299 46756 4355 46758
rect 4379 46756 4435 46758
rect 4459 46756 4515 46758
rect 4219 45722 4275 45724
rect 4299 45722 4355 45724
rect 4379 45722 4435 45724
rect 4459 45722 4515 45724
rect 4219 45670 4265 45722
rect 4265 45670 4275 45722
rect 4299 45670 4329 45722
rect 4329 45670 4341 45722
rect 4341 45670 4355 45722
rect 4379 45670 4393 45722
rect 4393 45670 4405 45722
rect 4405 45670 4435 45722
rect 4459 45670 4469 45722
rect 4469 45670 4515 45722
rect 4219 45668 4275 45670
rect 4299 45668 4355 45670
rect 4379 45668 4435 45670
rect 4459 45668 4515 45670
rect 3974 45056 4030 45112
rect 4219 44634 4275 44636
rect 4299 44634 4355 44636
rect 4379 44634 4435 44636
rect 4459 44634 4515 44636
rect 4219 44582 4265 44634
rect 4265 44582 4275 44634
rect 4299 44582 4329 44634
rect 4329 44582 4341 44634
rect 4341 44582 4355 44634
rect 4379 44582 4393 44634
rect 4393 44582 4405 44634
rect 4405 44582 4435 44634
rect 4459 44582 4469 44634
rect 4469 44582 4515 44634
rect 4219 44580 4275 44582
rect 4299 44580 4355 44582
rect 4379 44580 4435 44582
rect 4459 44580 4515 44582
rect 4219 43546 4275 43548
rect 4299 43546 4355 43548
rect 4379 43546 4435 43548
rect 4459 43546 4515 43548
rect 4219 43494 4265 43546
rect 4265 43494 4275 43546
rect 4299 43494 4329 43546
rect 4329 43494 4341 43546
rect 4341 43494 4355 43546
rect 4379 43494 4393 43546
rect 4393 43494 4405 43546
rect 4405 43494 4435 43546
rect 4459 43494 4469 43546
rect 4469 43494 4515 43546
rect 4219 43492 4275 43494
rect 4299 43492 4355 43494
rect 4379 43492 4435 43494
rect 4459 43492 4515 43494
rect 4219 42458 4275 42460
rect 4299 42458 4355 42460
rect 4379 42458 4435 42460
rect 4459 42458 4515 42460
rect 4219 42406 4265 42458
rect 4265 42406 4275 42458
rect 4299 42406 4329 42458
rect 4329 42406 4341 42458
rect 4341 42406 4355 42458
rect 4379 42406 4393 42458
rect 4393 42406 4405 42458
rect 4405 42406 4435 42458
rect 4459 42406 4469 42458
rect 4469 42406 4515 42458
rect 4219 42404 4275 42406
rect 4299 42404 4355 42406
rect 4379 42404 4435 42406
rect 4459 42404 4515 42406
rect 4066 41792 4122 41848
rect 4158 41540 4214 41576
rect 4158 41520 4160 41540
rect 4160 41520 4212 41540
rect 4212 41520 4214 41540
rect 4219 41370 4275 41372
rect 4299 41370 4355 41372
rect 4379 41370 4435 41372
rect 4459 41370 4515 41372
rect 4219 41318 4265 41370
rect 4265 41318 4275 41370
rect 4299 41318 4329 41370
rect 4329 41318 4341 41370
rect 4341 41318 4355 41370
rect 4379 41318 4393 41370
rect 4393 41318 4405 41370
rect 4405 41318 4435 41370
rect 4459 41318 4469 41370
rect 4469 41318 4515 41370
rect 4219 41316 4275 41318
rect 4299 41316 4355 41318
rect 4379 41316 4435 41318
rect 4459 41316 4515 41318
rect 4526 41112 4582 41168
rect 2588 23418 2644 23420
rect 2668 23418 2724 23420
rect 2748 23418 2804 23420
rect 2828 23418 2884 23420
rect 2588 23366 2634 23418
rect 2634 23366 2644 23418
rect 2668 23366 2698 23418
rect 2698 23366 2710 23418
rect 2710 23366 2724 23418
rect 2748 23366 2762 23418
rect 2762 23366 2774 23418
rect 2774 23366 2804 23418
rect 2828 23366 2838 23418
rect 2838 23366 2884 23418
rect 2588 23364 2644 23366
rect 2668 23364 2724 23366
rect 2748 23364 2804 23366
rect 2828 23364 2884 23366
rect 2588 22330 2644 22332
rect 2668 22330 2724 22332
rect 2748 22330 2804 22332
rect 2828 22330 2884 22332
rect 2588 22278 2634 22330
rect 2634 22278 2644 22330
rect 2668 22278 2698 22330
rect 2698 22278 2710 22330
rect 2710 22278 2724 22330
rect 2748 22278 2762 22330
rect 2762 22278 2774 22330
rect 2774 22278 2804 22330
rect 2828 22278 2838 22330
rect 2838 22278 2884 22330
rect 2588 22276 2644 22278
rect 2668 22276 2724 22278
rect 2748 22276 2804 22278
rect 2828 22276 2884 22278
rect 2588 21242 2644 21244
rect 2668 21242 2724 21244
rect 2748 21242 2804 21244
rect 2828 21242 2884 21244
rect 2588 21190 2634 21242
rect 2634 21190 2644 21242
rect 2668 21190 2698 21242
rect 2698 21190 2710 21242
rect 2710 21190 2724 21242
rect 2748 21190 2762 21242
rect 2762 21190 2774 21242
rect 2774 21190 2804 21242
rect 2828 21190 2838 21242
rect 2838 21190 2884 21242
rect 2588 21188 2644 21190
rect 2668 21188 2724 21190
rect 2748 21188 2804 21190
rect 2828 21188 2884 21190
rect 2588 20154 2644 20156
rect 2668 20154 2724 20156
rect 2748 20154 2804 20156
rect 2828 20154 2884 20156
rect 2588 20102 2634 20154
rect 2634 20102 2644 20154
rect 2668 20102 2698 20154
rect 2698 20102 2710 20154
rect 2710 20102 2724 20154
rect 2748 20102 2762 20154
rect 2762 20102 2774 20154
rect 2774 20102 2804 20154
rect 2828 20102 2838 20154
rect 2838 20102 2884 20154
rect 2588 20100 2644 20102
rect 2668 20100 2724 20102
rect 2748 20100 2804 20102
rect 2828 20100 2884 20102
rect 2588 19066 2644 19068
rect 2668 19066 2724 19068
rect 2748 19066 2804 19068
rect 2828 19066 2884 19068
rect 2588 19014 2634 19066
rect 2634 19014 2644 19066
rect 2668 19014 2698 19066
rect 2698 19014 2710 19066
rect 2710 19014 2724 19066
rect 2748 19014 2762 19066
rect 2762 19014 2774 19066
rect 2774 19014 2804 19066
rect 2828 19014 2838 19066
rect 2838 19014 2884 19066
rect 2588 19012 2644 19014
rect 2668 19012 2724 19014
rect 2748 19012 2804 19014
rect 2828 19012 2884 19014
rect 2588 17978 2644 17980
rect 2668 17978 2724 17980
rect 2748 17978 2804 17980
rect 2828 17978 2884 17980
rect 2588 17926 2634 17978
rect 2634 17926 2644 17978
rect 2668 17926 2698 17978
rect 2698 17926 2710 17978
rect 2710 17926 2724 17978
rect 2748 17926 2762 17978
rect 2762 17926 2774 17978
rect 2774 17926 2804 17978
rect 2828 17926 2838 17978
rect 2838 17926 2884 17978
rect 2588 17924 2644 17926
rect 2668 17924 2724 17926
rect 2748 17924 2804 17926
rect 2828 17924 2884 17926
rect 2588 16890 2644 16892
rect 2668 16890 2724 16892
rect 2748 16890 2804 16892
rect 2828 16890 2884 16892
rect 2588 16838 2634 16890
rect 2634 16838 2644 16890
rect 2668 16838 2698 16890
rect 2698 16838 2710 16890
rect 2710 16838 2724 16890
rect 2748 16838 2762 16890
rect 2762 16838 2774 16890
rect 2774 16838 2804 16890
rect 2828 16838 2838 16890
rect 2838 16838 2884 16890
rect 2588 16836 2644 16838
rect 2668 16836 2724 16838
rect 2748 16836 2804 16838
rect 2828 16836 2884 16838
rect 2588 15802 2644 15804
rect 2668 15802 2724 15804
rect 2748 15802 2804 15804
rect 2828 15802 2884 15804
rect 2588 15750 2634 15802
rect 2634 15750 2644 15802
rect 2668 15750 2698 15802
rect 2698 15750 2710 15802
rect 2710 15750 2724 15802
rect 2748 15750 2762 15802
rect 2762 15750 2774 15802
rect 2774 15750 2804 15802
rect 2828 15750 2838 15802
rect 2838 15750 2884 15802
rect 2588 15748 2644 15750
rect 2668 15748 2724 15750
rect 2748 15748 2804 15750
rect 2828 15748 2884 15750
rect 2588 14714 2644 14716
rect 2668 14714 2724 14716
rect 2748 14714 2804 14716
rect 2828 14714 2884 14716
rect 2588 14662 2634 14714
rect 2634 14662 2644 14714
rect 2668 14662 2698 14714
rect 2698 14662 2710 14714
rect 2710 14662 2724 14714
rect 2748 14662 2762 14714
rect 2762 14662 2774 14714
rect 2774 14662 2804 14714
rect 2828 14662 2838 14714
rect 2838 14662 2884 14714
rect 2588 14660 2644 14662
rect 2668 14660 2724 14662
rect 2748 14660 2804 14662
rect 2828 14660 2884 14662
rect 2588 13626 2644 13628
rect 2668 13626 2724 13628
rect 2748 13626 2804 13628
rect 2828 13626 2884 13628
rect 2588 13574 2634 13626
rect 2634 13574 2644 13626
rect 2668 13574 2698 13626
rect 2698 13574 2710 13626
rect 2710 13574 2724 13626
rect 2748 13574 2762 13626
rect 2762 13574 2774 13626
rect 2774 13574 2804 13626
rect 2828 13574 2838 13626
rect 2838 13574 2884 13626
rect 2588 13572 2644 13574
rect 2668 13572 2724 13574
rect 2748 13572 2804 13574
rect 2828 13572 2884 13574
rect 2588 12538 2644 12540
rect 2668 12538 2724 12540
rect 2748 12538 2804 12540
rect 2828 12538 2884 12540
rect 2588 12486 2634 12538
rect 2634 12486 2644 12538
rect 2668 12486 2698 12538
rect 2698 12486 2710 12538
rect 2710 12486 2724 12538
rect 2748 12486 2762 12538
rect 2762 12486 2774 12538
rect 2774 12486 2804 12538
rect 2828 12486 2838 12538
rect 2838 12486 2884 12538
rect 2588 12484 2644 12486
rect 2668 12484 2724 12486
rect 2748 12484 2804 12486
rect 2828 12484 2884 12486
rect 2588 11450 2644 11452
rect 2668 11450 2724 11452
rect 2748 11450 2804 11452
rect 2828 11450 2884 11452
rect 2588 11398 2634 11450
rect 2634 11398 2644 11450
rect 2668 11398 2698 11450
rect 2698 11398 2710 11450
rect 2710 11398 2724 11450
rect 2748 11398 2762 11450
rect 2762 11398 2774 11450
rect 2774 11398 2804 11450
rect 2828 11398 2838 11450
rect 2838 11398 2884 11450
rect 2588 11396 2644 11398
rect 2668 11396 2724 11398
rect 2748 11396 2804 11398
rect 2828 11396 2884 11398
rect 2588 10362 2644 10364
rect 2668 10362 2724 10364
rect 2748 10362 2804 10364
rect 2828 10362 2884 10364
rect 2588 10310 2634 10362
rect 2634 10310 2644 10362
rect 2668 10310 2698 10362
rect 2698 10310 2710 10362
rect 2710 10310 2724 10362
rect 2748 10310 2762 10362
rect 2762 10310 2774 10362
rect 2774 10310 2804 10362
rect 2828 10310 2838 10362
rect 2838 10310 2884 10362
rect 2588 10308 2644 10310
rect 2668 10308 2724 10310
rect 2748 10308 2804 10310
rect 2828 10308 2884 10310
rect 2588 9274 2644 9276
rect 2668 9274 2724 9276
rect 2748 9274 2804 9276
rect 2828 9274 2884 9276
rect 2588 9222 2634 9274
rect 2634 9222 2644 9274
rect 2668 9222 2698 9274
rect 2698 9222 2710 9274
rect 2710 9222 2724 9274
rect 2748 9222 2762 9274
rect 2762 9222 2774 9274
rect 2774 9222 2804 9274
rect 2828 9222 2838 9274
rect 2838 9222 2884 9274
rect 2588 9220 2644 9222
rect 2668 9220 2724 9222
rect 2748 9220 2804 9222
rect 2828 9220 2884 9222
rect 2318 9152 2374 9208
rect 2588 8186 2644 8188
rect 2668 8186 2724 8188
rect 2748 8186 2804 8188
rect 2828 8186 2884 8188
rect 2588 8134 2634 8186
rect 2634 8134 2644 8186
rect 2668 8134 2698 8186
rect 2698 8134 2710 8186
rect 2710 8134 2724 8186
rect 2748 8134 2762 8186
rect 2762 8134 2774 8186
rect 2774 8134 2804 8186
rect 2828 8134 2838 8186
rect 2838 8134 2884 8186
rect 2588 8132 2644 8134
rect 2668 8132 2724 8134
rect 2748 8132 2804 8134
rect 2828 8132 2884 8134
rect 1490 5208 1546 5264
rect 1490 4664 1546 4720
rect 1490 4120 1546 4176
rect 2042 6976 2098 7032
rect 1490 3032 1546 3088
rect 1398 2488 1454 2544
rect 2588 7098 2644 7100
rect 2668 7098 2724 7100
rect 2748 7098 2804 7100
rect 2828 7098 2884 7100
rect 2588 7046 2634 7098
rect 2634 7046 2644 7098
rect 2668 7046 2698 7098
rect 2698 7046 2710 7098
rect 2710 7046 2724 7098
rect 2748 7046 2762 7098
rect 2762 7046 2774 7098
rect 2774 7046 2804 7098
rect 2828 7046 2838 7098
rect 2838 7046 2884 7098
rect 2588 7044 2644 7046
rect 2668 7044 2724 7046
rect 2748 7044 2804 7046
rect 2828 7044 2884 7046
rect 4219 40282 4275 40284
rect 4299 40282 4355 40284
rect 4379 40282 4435 40284
rect 4459 40282 4515 40284
rect 4219 40230 4265 40282
rect 4265 40230 4275 40282
rect 4299 40230 4329 40282
rect 4329 40230 4341 40282
rect 4341 40230 4355 40282
rect 4379 40230 4393 40282
rect 4393 40230 4405 40282
rect 4405 40230 4435 40282
rect 4459 40230 4469 40282
rect 4469 40230 4515 40282
rect 4219 40228 4275 40230
rect 4299 40228 4355 40230
rect 4379 40228 4435 40230
rect 4459 40228 4515 40230
rect 4219 39194 4275 39196
rect 4299 39194 4355 39196
rect 4379 39194 4435 39196
rect 4459 39194 4515 39196
rect 4219 39142 4265 39194
rect 4265 39142 4275 39194
rect 4299 39142 4329 39194
rect 4329 39142 4341 39194
rect 4341 39142 4355 39194
rect 4379 39142 4393 39194
rect 4393 39142 4405 39194
rect 4405 39142 4435 39194
rect 4459 39142 4469 39194
rect 4469 39142 4515 39194
rect 4219 39140 4275 39142
rect 4299 39140 4355 39142
rect 4379 39140 4435 39142
rect 4459 39140 4515 39142
rect 4219 38106 4275 38108
rect 4299 38106 4355 38108
rect 4379 38106 4435 38108
rect 4459 38106 4515 38108
rect 4219 38054 4265 38106
rect 4265 38054 4275 38106
rect 4299 38054 4329 38106
rect 4329 38054 4341 38106
rect 4341 38054 4355 38106
rect 4379 38054 4393 38106
rect 4393 38054 4405 38106
rect 4405 38054 4435 38106
rect 4459 38054 4469 38106
rect 4469 38054 4515 38106
rect 4219 38052 4275 38054
rect 4299 38052 4355 38054
rect 4379 38052 4435 38054
rect 4459 38052 4515 38054
rect 4219 37018 4275 37020
rect 4299 37018 4355 37020
rect 4379 37018 4435 37020
rect 4459 37018 4515 37020
rect 4219 36966 4265 37018
rect 4265 36966 4275 37018
rect 4299 36966 4329 37018
rect 4329 36966 4341 37018
rect 4341 36966 4355 37018
rect 4379 36966 4393 37018
rect 4393 36966 4405 37018
rect 4405 36966 4435 37018
rect 4459 36966 4469 37018
rect 4469 36966 4515 37018
rect 4219 36964 4275 36966
rect 4299 36964 4355 36966
rect 4379 36964 4435 36966
rect 4459 36964 4515 36966
rect 4219 35930 4275 35932
rect 4299 35930 4355 35932
rect 4379 35930 4435 35932
rect 4459 35930 4515 35932
rect 4219 35878 4265 35930
rect 4265 35878 4275 35930
rect 4299 35878 4329 35930
rect 4329 35878 4341 35930
rect 4341 35878 4355 35930
rect 4379 35878 4393 35930
rect 4393 35878 4405 35930
rect 4405 35878 4435 35930
rect 4459 35878 4469 35930
rect 4469 35878 4515 35930
rect 4219 35876 4275 35878
rect 4299 35876 4355 35878
rect 4379 35876 4435 35878
rect 4459 35876 4515 35878
rect 4219 34842 4275 34844
rect 4299 34842 4355 34844
rect 4379 34842 4435 34844
rect 4459 34842 4515 34844
rect 4219 34790 4265 34842
rect 4265 34790 4275 34842
rect 4299 34790 4329 34842
rect 4329 34790 4341 34842
rect 4341 34790 4355 34842
rect 4379 34790 4393 34842
rect 4393 34790 4405 34842
rect 4405 34790 4435 34842
rect 4459 34790 4469 34842
rect 4469 34790 4515 34842
rect 4219 34788 4275 34790
rect 4299 34788 4355 34790
rect 4379 34788 4435 34790
rect 4459 34788 4515 34790
rect 4618 34312 4674 34368
rect 4219 33754 4275 33756
rect 4299 33754 4355 33756
rect 4379 33754 4435 33756
rect 4459 33754 4515 33756
rect 4219 33702 4265 33754
rect 4265 33702 4275 33754
rect 4299 33702 4329 33754
rect 4329 33702 4341 33754
rect 4341 33702 4355 33754
rect 4379 33702 4393 33754
rect 4393 33702 4405 33754
rect 4405 33702 4435 33754
rect 4459 33702 4469 33754
rect 4469 33702 4515 33754
rect 4219 33700 4275 33702
rect 4299 33700 4355 33702
rect 4379 33700 4435 33702
rect 4459 33700 4515 33702
rect 4219 32666 4275 32668
rect 4299 32666 4355 32668
rect 4379 32666 4435 32668
rect 4459 32666 4515 32668
rect 4219 32614 4265 32666
rect 4265 32614 4275 32666
rect 4299 32614 4329 32666
rect 4329 32614 4341 32666
rect 4341 32614 4355 32666
rect 4379 32614 4393 32666
rect 4393 32614 4405 32666
rect 4405 32614 4435 32666
rect 4459 32614 4469 32666
rect 4469 32614 4515 32666
rect 4219 32612 4275 32614
rect 4299 32612 4355 32614
rect 4379 32612 4435 32614
rect 4459 32612 4515 32614
rect 4219 31578 4275 31580
rect 4299 31578 4355 31580
rect 4379 31578 4435 31580
rect 4459 31578 4515 31580
rect 4219 31526 4265 31578
rect 4265 31526 4275 31578
rect 4299 31526 4329 31578
rect 4329 31526 4341 31578
rect 4341 31526 4355 31578
rect 4379 31526 4393 31578
rect 4393 31526 4405 31578
rect 4405 31526 4435 31578
rect 4459 31526 4469 31578
rect 4469 31526 4515 31578
rect 4219 31524 4275 31526
rect 4299 31524 4355 31526
rect 4379 31524 4435 31526
rect 4459 31524 4515 31526
rect 4219 30490 4275 30492
rect 4299 30490 4355 30492
rect 4379 30490 4435 30492
rect 4459 30490 4515 30492
rect 4219 30438 4265 30490
rect 4265 30438 4275 30490
rect 4299 30438 4329 30490
rect 4329 30438 4341 30490
rect 4341 30438 4355 30490
rect 4379 30438 4393 30490
rect 4393 30438 4405 30490
rect 4405 30438 4435 30490
rect 4459 30438 4469 30490
rect 4469 30438 4515 30490
rect 4219 30436 4275 30438
rect 4299 30436 4355 30438
rect 4379 30436 4435 30438
rect 4459 30436 4515 30438
rect 4219 29402 4275 29404
rect 4299 29402 4355 29404
rect 4379 29402 4435 29404
rect 4459 29402 4515 29404
rect 4219 29350 4265 29402
rect 4265 29350 4275 29402
rect 4299 29350 4329 29402
rect 4329 29350 4341 29402
rect 4341 29350 4355 29402
rect 4379 29350 4393 29402
rect 4393 29350 4405 29402
rect 4405 29350 4435 29402
rect 4459 29350 4469 29402
rect 4469 29350 4515 29402
rect 4219 29348 4275 29350
rect 4299 29348 4355 29350
rect 4379 29348 4435 29350
rect 4459 29348 4515 29350
rect 4219 28314 4275 28316
rect 4299 28314 4355 28316
rect 4379 28314 4435 28316
rect 4459 28314 4515 28316
rect 4219 28262 4265 28314
rect 4265 28262 4275 28314
rect 4299 28262 4329 28314
rect 4329 28262 4341 28314
rect 4341 28262 4355 28314
rect 4379 28262 4393 28314
rect 4393 28262 4405 28314
rect 4405 28262 4435 28314
rect 4459 28262 4469 28314
rect 4469 28262 4515 28314
rect 4219 28260 4275 28262
rect 4299 28260 4355 28262
rect 4379 28260 4435 28262
rect 4459 28260 4515 28262
rect 4219 27226 4275 27228
rect 4299 27226 4355 27228
rect 4379 27226 4435 27228
rect 4459 27226 4515 27228
rect 4219 27174 4265 27226
rect 4265 27174 4275 27226
rect 4299 27174 4329 27226
rect 4329 27174 4341 27226
rect 4341 27174 4355 27226
rect 4379 27174 4393 27226
rect 4393 27174 4405 27226
rect 4405 27174 4435 27226
rect 4459 27174 4469 27226
rect 4469 27174 4515 27226
rect 4219 27172 4275 27174
rect 4299 27172 4355 27174
rect 4379 27172 4435 27174
rect 4459 27172 4515 27174
rect 4219 26138 4275 26140
rect 4299 26138 4355 26140
rect 4379 26138 4435 26140
rect 4459 26138 4515 26140
rect 4219 26086 4265 26138
rect 4265 26086 4275 26138
rect 4299 26086 4329 26138
rect 4329 26086 4341 26138
rect 4341 26086 4355 26138
rect 4379 26086 4393 26138
rect 4393 26086 4405 26138
rect 4405 26086 4435 26138
rect 4459 26086 4469 26138
rect 4469 26086 4515 26138
rect 4219 26084 4275 26086
rect 4299 26084 4355 26086
rect 4379 26084 4435 26086
rect 4459 26084 4515 26086
rect 4219 25050 4275 25052
rect 4299 25050 4355 25052
rect 4379 25050 4435 25052
rect 4459 25050 4515 25052
rect 4219 24998 4265 25050
rect 4265 24998 4275 25050
rect 4299 24998 4329 25050
rect 4329 24998 4341 25050
rect 4341 24998 4355 25050
rect 4379 24998 4393 25050
rect 4393 24998 4405 25050
rect 4405 24998 4435 25050
rect 4459 24998 4469 25050
rect 4469 24998 4515 25050
rect 4219 24996 4275 24998
rect 4299 24996 4355 24998
rect 4379 24996 4435 24998
rect 4459 24996 4515 24998
rect 4219 23962 4275 23964
rect 4299 23962 4355 23964
rect 4379 23962 4435 23964
rect 4459 23962 4515 23964
rect 4219 23910 4265 23962
rect 4265 23910 4275 23962
rect 4299 23910 4329 23962
rect 4329 23910 4341 23962
rect 4341 23910 4355 23962
rect 4379 23910 4393 23962
rect 4393 23910 4405 23962
rect 4405 23910 4435 23962
rect 4459 23910 4469 23962
rect 4469 23910 4515 23962
rect 4219 23908 4275 23910
rect 4299 23908 4355 23910
rect 4379 23908 4435 23910
rect 4459 23908 4515 23910
rect 4219 22874 4275 22876
rect 4299 22874 4355 22876
rect 4379 22874 4435 22876
rect 4459 22874 4515 22876
rect 4219 22822 4265 22874
rect 4265 22822 4275 22874
rect 4299 22822 4329 22874
rect 4329 22822 4341 22874
rect 4341 22822 4355 22874
rect 4379 22822 4393 22874
rect 4393 22822 4405 22874
rect 4405 22822 4435 22874
rect 4459 22822 4469 22874
rect 4469 22822 4515 22874
rect 4219 22820 4275 22822
rect 4299 22820 4355 22822
rect 4379 22820 4435 22822
rect 4459 22820 4515 22822
rect 4219 21786 4275 21788
rect 4299 21786 4355 21788
rect 4379 21786 4435 21788
rect 4459 21786 4515 21788
rect 4219 21734 4265 21786
rect 4265 21734 4275 21786
rect 4299 21734 4329 21786
rect 4329 21734 4341 21786
rect 4341 21734 4355 21786
rect 4379 21734 4393 21786
rect 4393 21734 4405 21786
rect 4405 21734 4435 21786
rect 4459 21734 4469 21786
rect 4469 21734 4515 21786
rect 4219 21732 4275 21734
rect 4299 21732 4355 21734
rect 4379 21732 4435 21734
rect 4459 21732 4515 21734
rect 4219 20698 4275 20700
rect 4299 20698 4355 20700
rect 4379 20698 4435 20700
rect 4459 20698 4515 20700
rect 4219 20646 4265 20698
rect 4265 20646 4275 20698
rect 4299 20646 4329 20698
rect 4329 20646 4341 20698
rect 4341 20646 4355 20698
rect 4379 20646 4393 20698
rect 4393 20646 4405 20698
rect 4405 20646 4435 20698
rect 4459 20646 4469 20698
rect 4469 20646 4515 20698
rect 4219 20644 4275 20646
rect 4299 20644 4355 20646
rect 4379 20644 4435 20646
rect 4459 20644 4515 20646
rect 4219 19610 4275 19612
rect 4299 19610 4355 19612
rect 4379 19610 4435 19612
rect 4459 19610 4515 19612
rect 4219 19558 4265 19610
rect 4265 19558 4275 19610
rect 4299 19558 4329 19610
rect 4329 19558 4341 19610
rect 4341 19558 4355 19610
rect 4379 19558 4393 19610
rect 4393 19558 4405 19610
rect 4405 19558 4435 19610
rect 4459 19558 4469 19610
rect 4469 19558 4515 19610
rect 4219 19556 4275 19558
rect 4299 19556 4355 19558
rect 4379 19556 4435 19558
rect 4459 19556 4515 19558
rect 4219 18522 4275 18524
rect 4299 18522 4355 18524
rect 4379 18522 4435 18524
rect 4459 18522 4515 18524
rect 4219 18470 4265 18522
rect 4265 18470 4275 18522
rect 4299 18470 4329 18522
rect 4329 18470 4341 18522
rect 4341 18470 4355 18522
rect 4379 18470 4393 18522
rect 4393 18470 4405 18522
rect 4405 18470 4435 18522
rect 4459 18470 4469 18522
rect 4469 18470 4515 18522
rect 4219 18468 4275 18470
rect 4299 18468 4355 18470
rect 4379 18468 4435 18470
rect 4459 18468 4515 18470
rect 4219 17434 4275 17436
rect 4299 17434 4355 17436
rect 4379 17434 4435 17436
rect 4459 17434 4515 17436
rect 4219 17382 4265 17434
rect 4265 17382 4275 17434
rect 4299 17382 4329 17434
rect 4329 17382 4341 17434
rect 4341 17382 4355 17434
rect 4379 17382 4393 17434
rect 4393 17382 4405 17434
rect 4405 17382 4435 17434
rect 4459 17382 4469 17434
rect 4469 17382 4515 17434
rect 4219 17380 4275 17382
rect 4299 17380 4355 17382
rect 4379 17380 4435 17382
rect 4459 17380 4515 17382
rect 4219 16346 4275 16348
rect 4299 16346 4355 16348
rect 4379 16346 4435 16348
rect 4459 16346 4515 16348
rect 4219 16294 4265 16346
rect 4265 16294 4275 16346
rect 4299 16294 4329 16346
rect 4329 16294 4341 16346
rect 4341 16294 4355 16346
rect 4379 16294 4393 16346
rect 4393 16294 4405 16346
rect 4405 16294 4435 16346
rect 4459 16294 4469 16346
rect 4469 16294 4515 16346
rect 4219 16292 4275 16294
rect 4299 16292 4355 16294
rect 4379 16292 4435 16294
rect 4459 16292 4515 16294
rect 4219 15258 4275 15260
rect 4299 15258 4355 15260
rect 4379 15258 4435 15260
rect 4459 15258 4515 15260
rect 4219 15206 4265 15258
rect 4265 15206 4275 15258
rect 4299 15206 4329 15258
rect 4329 15206 4341 15258
rect 4341 15206 4355 15258
rect 4379 15206 4393 15258
rect 4393 15206 4405 15258
rect 4405 15206 4435 15258
rect 4459 15206 4469 15258
rect 4469 15206 4515 15258
rect 4219 15204 4275 15206
rect 4299 15204 4355 15206
rect 4379 15204 4435 15206
rect 4459 15204 4515 15206
rect 4219 14170 4275 14172
rect 4299 14170 4355 14172
rect 4379 14170 4435 14172
rect 4459 14170 4515 14172
rect 4219 14118 4265 14170
rect 4265 14118 4275 14170
rect 4299 14118 4329 14170
rect 4329 14118 4341 14170
rect 4341 14118 4355 14170
rect 4379 14118 4393 14170
rect 4393 14118 4405 14170
rect 4405 14118 4435 14170
rect 4459 14118 4469 14170
rect 4469 14118 4515 14170
rect 4219 14116 4275 14118
rect 4299 14116 4355 14118
rect 4379 14116 4435 14118
rect 4459 14116 4515 14118
rect 4219 13082 4275 13084
rect 4299 13082 4355 13084
rect 4379 13082 4435 13084
rect 4459 13082 4515 13084
rect 4219 13030 4265 13082
rect 4265 13030 4275 13082
rect 4299 13030 4329 13082
rect 4329 13030 4341 13082
rect 4341 13030 4355 13082
rect 4379 13030 4393 13082
rect 4393 13030 4405 13082
rect 4405 13030 4435 13082
rect 4459 13030 4469 13082
rect 4469 13030 4515 13082
rect 4219 13028 4275 13030
rect 4299 13028 4355 13030
rect 4379 13028 4435 13030
rect 4459 13028 4515 13030
rect 2588 6010 2644 6012
rect 2668 6010 2724 6012
rect 2748 6010 2804 6012
rect 2828 6010 2884 6012
rect 2588 5958 2634 6010
rect 2634 5958 2644 6010
rect 2668 5958 2698 6010
rect 2698 5958 2710 6010
rect 2710 5958 2724 6010
rect 2748 5958 2762 6010
rect 2762 5958 2774 6010
rect 2774 5958 2804 6010
rect 2828 5958 2838 6010
rect 2838 5958 2884 6010
rect 2588 5956 2644 5958
rect 2668 5956 2724 5958
rect 2748 5956 2804 5958
rect 2828 5956 2884 5958
rect 2588 4922 2644 4924
rect 2668 4922 2724 4924
rect 2748 4922 2804 4924
rect 2828 4922 2884 4924
rect 2588 4870 2634 4922
rect 2634 4870 2644 4922
rect 2668 4870 2698 4922
rect 2698 4870 2710 4922
rect 2710 4870 2724 4922
rect 2748 4870 2762 4922
rect 2762 4870 2774 4922
rect 2774 4870 2804 4922
rect 2828 4870 2838 4922
rect 2838 4870 2884 4922
rect 2588 4868 2644 4870
rect 2668 4868 2724 4870
rect 2748 4868 2804 4870
rect 2828 4868 2884 4870
rect 2588 3834 2644 3836
rect 2668 3834 2724 3836
rect 2748 3834 2804 3836
rect 2828 3834 2884 3836
rect 2588 3782 2634 3834
rect 2634 3782 2644 3834
rect 2668 3782 2698 3834
rect 2698 3782 2710 3834
rect 2710 3782 2724 3834
rect 2748 3782 2762 3834
rect 2762 3782 2774 3834
rect 2774 3782 2804 3834
rect 2828 3782 2838 3834
rect 2838 3782 2884 3834
rect 2588 3780 2644 3782
rect 2668 3780 2724 3782
rect 2748 3780 2804 3782
rect 2828 3780 2884 3782
rect 2318 3576 2374 3632
rect 4219 11994 4275 11996
rect 4299 11994 4355 11996
rect 4379 11994 4435 11996
rect 4459 11994 4515 11996
rect 4219 11942 4265 11994
rect 4265 11942 4275 11994
rect 4299 11942 4329 11994
rect 4329 11942 4341 11994
rect 4341 11942 4355 11994
rect 4379 11942 4393 11994
rect 4393 11942 4405 11994
rect 4405 11942 4435 11994
rect 4459 11942 4469 11994
rect 4469 11942 4515 11994
rect 4219 11940 4275 11942
rect 4299 11940 4355 11942
rect 4379 11940 4435 11942
rect 4459 11940 4515 11942
rect 4219 10906 4275 10908
rect 4299 10906 4355 10908
rect 4379 10906 4435 10908
rect 4459 10906 4515 10908
rect 4219 10854 4265 10906
rect 4265 10854 4275 10906
rect 4299 10854 4329 10906
rect 4329 10854 4341 10906
rect 4341 10854 4355 10906
rect 4379 10854 4393 10906
rect 4393 10854 4405 10906
rect 4405 10854 4435 10906
rect 4459 10854 4469 10906
rect 4469 10854 4515 10906
rect 4219 10852 4275 10854
rect 4299 10852 4355 10854
rect 4379 10852 4435 10854
rect 4459 10852 4515 10854
rect 4219 9818 4275 9820
rect 4299 9818 4355 9820
rect 4379 9818 4435 9820
rect 4459 9818 4515 9820
rect 4219 9766 4265 9818
rect 4265 9766 4275 9818
rect 4299 9766 4329 9818
rect 4329 9766 4341 9818
rect 4341 9766 4355 9818
rect 4379 9766 4393 9818
rect 4393 9766 4405 9818
rect 4405 9766 4435 9818
rect 4459 9766 4469 9818
rect 4469 9766 4515 9818
rect 4219 9764 4275 9766
rect 4299 9764 4355 9766
rect 4379 9764 4435 9766
rect 4459 9764 4515 9766
rect 4219 8730 4275 8732
rect 4299 8730 4355 8732
rect 4379 8730 4435 8732
rect 4459 8730 4515 8732
rect 4219 8678 4265 8730
rect 4265 8678 4275 8730
rect 4299 8678 4329 8730
rect 4329 8678 4341 8730
rect 4341 8678 4355 8730
rect 4379 8678 4393 8730
rect 4393 8678 4405 8730
rect 4405 8678 4435 8730
rect 4459 8678 4469 8730
rect 4469 8678 4515 8730
rect 4219 8676 4275 8678
rect 4299 8676 4355 8678
rect 4379 8676 4435 8678
rect 4459 8676 4515 8678
rect 4219 7642 4275 7644
rect 4299 7642 4355 7644
rect 4379 7642 4435 7644
rect 4459 7642 4515 7644
rect 4219 7590 4265 7642
rect 4265 7590 4275 7642
rect 4299 7590 4329 7642
rect 4329 7590 4341 7642
rect 4341 7590 4355 7642
rect 4379 7590 4393 7642
rect 4393 7590 4405 7642
rect 4405 7590 4435 7642
rect 4459 7590 4469 7642
rect 4469 7590 4515 7642
rect 4219 7588 4275 7590
rect 4299 7588 4355 7590
rect 4379 7588 4435 7590
rect 4459 7588 4515 7590
rect 4219 6554 4275 6556
rect 4299 6554 4355 6556
rect 4379 6554 4435 6556
rect 4459 6554 4515 6556
rect 4219 6502 4265 6554
rect 4265 6502 4275 6554
rect 4299 6502 4329 6554
rect 4329 6502 4341 6554
rect 4341 6502 4355 6554
rect 4379 6502 4393 6554
rect 4393 6502 4405 6554
rect 4405 6502 4435 6554
rect 4459 6502 4469 6554
rect 4469 6502 4515 6554
rect 4219 6500 4275 6502
rect 4299 6500 4355 6502
rect 4379 6500 4435 6502
rect 4459 6500 4515 6502
rect 5078 39888 5134 39944
rect 5262 39344 5318 39400
rect 5354 35808 5410 35864
rect 5851 73466 5907 73468
rect 5931 73466 5987 73468
rect 6011 73466 6067 73468
rect 6091 73466 6147 73468
rect 5851 73414 5897 73466
rect 5897 73414 5907 73466
rect 5931 73414 5961 73466
rect 5961 73414 5973 73466
rect 5973 73414 5987 73466
rect 6011 73414 6025 73466
rect 6025 73414 6037 73466
rect 6037 73414 6067 73466
rect 6091 73414 6101 73466
rect 6101 73414 6147 73466
rect 5851 73412 5907 73414
rect 5931 73412 5987 73414
rect 6011 73412 6067 73414
rect 6091 73412 6147 73414
rect 5078 35400 5134 35456
rect 5851 72378 5907 72380
rect 5931 72378 5987 72380
rect 6011 72378 6067 72380
rect 6091 72378 6147 72380
rect 5851 72326 5897 72378
rect 5897 72326 5907 72378
rect 5931 72326 5961 72378
rect 5961 72326 5973 72378
rect 5973 72326 5987 72378
rect 6011 72326 6025 72378
rect 6025 72326 6037 72378
rect 6037 72326 6067 72378
rect 6091 72326 6101 72378
rect 6101 72326 6147 72378
rect 5851 72324 5907 72326
rect 5931 72324 5987 72326
rect 6011 72324 6067 72326
rect 6091 72324 6147 72326
rect 5851 71290 5907 71292
rect 5931 71290 5987 71292
rect 6011 71290 6067 71292
rect 6091 71290 6147 71292
rect 5851 71238 5897 71290
rect 5897 71238 5907 71290
rect 5931 71238 5961 71290
rect 5961 71238 5973 71290
rect 5973 71238 5987 71290
rect 6011 71238 6025 71290
rect 6025 71238 6037 71290
rect 6037 71238 6067 71290
rect 6091 71238 6101 71290
rect 6101 71238 6147 71290
rect 5851 71236 5907 71238
rect 5931 71236 5987 71238
rect 6011 71236 6067 71238
rect 6091 71236 6147 71238
rect 5851 70202 5907 70204
rect 5931 70202 5987 70204
rect 6011 70202 6067 70204
rect 6091 70202 6147 70204
rect 5851 70150 5897 70202
rect 5897 70150 5907 70202
rect 5931 70150 5961 70202
rect 5961 70150 5973 70202
rect 5973 70150 5987 70202
rect 6011 70150 6025 70202
rect 6025 70150 6037 70202
rect 6037 70150 6067 70202
rect 6091 70150 6101 70202
rect 6101 70150 6147 70202
rect 5851 70148 5907 70150
rect 5931 70148 5987 70150
rect 6011 70148 6067 70150
rect 6091 70148 6147 70150
rect 5851 69114 5907 69116
rect 5931 69114 5987 69116
rect 6011 69114 6067 69116
rect 6091 69114 6147 69116
rect 5851 69062 5897 69114
rect 5897 69062 5907 69114
rect 5931 69062 5961 69114
rect 5961 69062 5973 69114
rect 5973 69062 5987 69114
rect 6011 69062 6025 69114
rect 6025 69062 6037 69114
rect 6037 69062 6067 69114
rect 6091 69062 6101 69114
rect 6101 69062 6147 69114
rect 5851 69060 5907 69062
rect 5931 69060 5987 69062
rect 6011 69060 6067 69062
rect 6091 69060 6147 69062
rect 5851 68026 5907 68028
rect 5931 68026 5987 68028
rect 6011 68026 6067 68028
rect 6091 68026 6147 68028
rect 5851 67974 5897 68026
rect 5897 67974 5907 68026
rect 5931 67974 5961 68026
rect 5961 67974 5973 68026
rect 5973 67974 5987 68026
rect 6011 67974 6025 68026
rect 6025 67974 6037 68026
rect 6037 67974 6067 68026
rect 6091 67974 6101 68026
rect 6101 67974 6147 68026
rect 5851 67972 5907 67974
rect 5931 67972 5987 67974
rect 6011 67972 6067 67974
rect 6091 67972 6147 67974
rect 5851 66938 5907 66940
rect 5931 66938 5987 66940
rect 6011 66938 6067 66940
rect 6091 66938 6147 66940
rect 5851 66886 5897 66938
rect 5897 66886 5907 66938
rect 5931 66886 5961 66938
rect 5961 66886 5973 66938
rect 5973 66886 5987 66938
rect 6011 66886 6025 66938
rect 6025 66886 6037 66938
rect 6037 66886 6067 66938
rect 6091 66886 6101 66938
rect 6101 66886 6147 66938
rect 5851 66884 5907 66886
rect 5931 66884 5987 66886
rect 6011 66884 6067 66886
rect 6091 66884 6147 66886
rect 5851 65850 5907 65852
rect 5931 65850 5987 65852
rect 6011 65850 6067 65852
rect 6091 65850 6147 65852
rect 5851 65798 5897 65850
rect 5897 65798 5907 65850
rect 5931 65798 5961 65850
rect 5961 65798 5973 65850
rect 5973 65798 5987 65850
rect 6011 65798 6025 65850
rect 6025 65798 6037 65850
rect 6037 65798 6067 65850
rect 6091 65798 6101 65850
rect 6101 65798 6147 65850
rect 5851 65796 5907 65798
rect 5931 65796 5987 65798
rect 6011 65796 6067 65798
rect 6091 65796 6147 65798
rect 5851 64762 5907 64764
rect 5931 64762 5987 64764
rect 6011 64762 6067 64764
rect 6091 64762 6147 64764
rect 5851 64710 5897 64762
rect 5897 64710 5907 64762
rect 5931 64710 5961 64762
rect 5961 64710 5973 64762
rect 5973 64710 5987 64762
rect 6011 64710 6025 64762
rect 6025 64710 6037 64762
rect 6037 64710 6067 64762
rect 6091 64710 6101 64762
rect 6101 64710 6147 64762
rect 5851 64708 5907 64710
rect 5931 64708 5987 64710
rect 6011 64708 6067 64710
rect 6091 64708 6147 64710
rect 5851 63674 5907 63676
rect 5931 63674 5987 63676
rect 6011 63674 6067 63676
rect 6091 63674 6147 63676
rect 5851 63622 5897 63674
rect 5897 63622 5907 63674
rect 5931 63622 5961 63674
rect 5961 63622 5973 63674
rect 5973 63622 5987 63674
rect 6011 63622 6025 63674
rect 6025 63622 6037 63674
rect 6037 63622 6067 63674
rect 6091 63622 6101 63674
rect 6101 63622 6147 63674
rect 5851 63620 5907 63622
rect 5931 63620 5987 63622
rect 6011 63620 6067 63622
rect 6091 63620 6147 63622
rect 5851 62586 5907 62588
rect 5931 62586 5987 62588
rect 6011 62586 6067 62588
rect 6091 62586 6147 62588
rect 5851 62534 5897 62586
rect 5897 62534 5907 62586
rect 5931 62534 5961 62586
rect 5961 62534 5973 62586
rect 5973 62534 5987 62586
rect 6011 62534 6025 62586
rect 6025 62534 6037 62586
rect 6037 62534 6067 62586
rect 6091 62534 6101 62586
rect 6101 62534 6147 62586
rect 5851 62532 5907 62534
rect 5931 62532 5987 62534
rect 6011 62532 6067 62534
rect 6091 62532 6147 62534
rect 5851 61498 5907 61500
rect 5931 61498 5987 61500
rect 6011 61498 6067 61500
rect 6091 61498 6147 61500
rect 5851 61446 5897 61498
rect 5897 61446 5907 61498
rect 5931 61446 5961 61498
rect 5961 61446 5973 61498
rect 5973 61446 5987 61498
rect 6011 61446 6025 61498
rect 6025 61446 6037 61498
rect 6037 61446 6067 61498
rect 6091 61446 6101 61498
rect 6101 61446 6147 61498
rect 5851 61444 5907 61446
rect 5931 61444 5987 61446
rect 6011 61444 6067 61446
rect 6091 61444 6147 61446
rect 5851 60410 5907 60412
rect 5931 60410 5987 60412
rect 6011 60410 6067 60412
rect 6091 60410 6147 60412
rect 5851 60358 5897 60410
rect 5897 60358 5907 60410
rect 5931 60358 5961 60410
rect 5961 60358 5973 60410
rect 5973 60358 5987 60410
rect 6011 60358 6025 60410
rect 6025 60358 6037 60410
rect 6037 60358 6067 60410
rect 6091 60358 6101 60410
rect 6101 60358 6147 60410
rect 5851 60356 5907 60358
rect 5931 60356 5987 60358
rect 6011 60356 6067 60358
rect 6091 60356 6147 60358
rect 5851 59322 5907 59324
rect 5931 59322 5987 59324
rect 6011 59322 6067 59324
rect 6091 59322 6147 59324
rect 5851 59270 5897 59322
rect 5897 59270 5907 59322
rect 5931 59270 5961 59322
rect 5961 59270 5973 59322
rect 5973 59270 5987 59322
rect 6011 59270 6025 59322
rect 6025 59270 6037 59322
rect 6037 59270 6067 59322
rect 6091 59270 6101 59322
rect 6101 59270 6147 59322
rect 5851 59268 5907 59270
rect 5931 59268 5987 59270
rect 6011 59268 6067 59270
rect 6091 59268 6147 59270
rect 5851 58234 5907 58236
rect 5931 58234 5987 58236
rect 6011 58234 6067 58236
rect 6091 58234 6147 58236
rect 5851 58182 5897 58234
rect 5897 58182 5907 58234
rect 5931 58182 5961 58234
rect 5961 58182 5973 58234
rect 5973 58182 5987 58234
rect 6011 58182 6025 58234
rect 6025 58182 6037 58234
rect 6037 58182 6067 58234
rect 6091 58182 6101 58234
rect 6101 58182 6147 58234
rect 5851 58180 5907 58182
rect 5931 58180 5987 58182
rect 6011 58180 6067 58182
rect 6091 58180 6147 58182
rect 5851 57146 5907 57148
rect 5931 57146 5987 57148
rect 6011 57146 6067 57148
rect 6091 57146 6147 57148
rect 5851 57094 5897 57146
rect 5897 57094 5907 57146
rect 5931 57094 5961 57146
rect 5961 57094 5973 57146
rect 5973 57094 5987 57146
rect 6011 57094 6025 57146
rect 6025 57094 6037 57146
rect 6037 57094 6067 57146
rect 6091 57094 6101 57146
rect 6101 57094 6147 57146
rect 5851 57092 5907 57094
rect 5931 57092 5987 57094
rect 6011 57092 6067 57094
rect 6091 57092 6147 57094
rect 5814 56208 5870 56264
rect 5851 56058 5907 56060
rect 5931 56058 5987 56060
rect 6011 56058 6067 56060
rect 6091 56058 6147 56060
rect 5851 56006 5897 56058
rect 5897 56006 5907 56058
rect 5931 56006 5961 56058
rect 5961 56006 5973 56058
rect 5973 56006 5987 56058
rect 6011 56006 6025 56058
rect 6025 56006 6037 56058
rect 6037 56006 6067 56058
rect 6091 56006 6101 56058
rect 6101 56006 6147 56058
rect 5851 56004 5907 56006
rect 5931 56004 5987 56006
rect 6011 56004 6067 56006
rect 6091 56004 6147 56006
rect 5851 54970 5907 54972
rect 5931 54970 5987 54972
rect 6011 54970 6067 54972
rect 6091 54970 6147 54972
rect 5851 54918 5897 54970
rect 5897 54918 5907 54970
rect 5931 54918 5961 54970
rect 5961 54918 5973 54970
rect 5973 54918 5987 54970
rect 6011 54918 6025 54970
rect 6025 54918 6037 54970
rect 6037 54918 6067 54970
rect 6091 54918 6101 54970
rect 6101 54918 6147 54970
rect 5851 54916 5907 54918
rect 5931 54916 5987 54918
rect 6011 54916 6067 54918
rect 6091 54916 6147 54918
rect 5851 53882 5907 53884
rect 5931 53882 5987 53884
rect 6011 53882 6067 53884
rect 6091 53882 6147 53884
rect 5851 53830 5897 53882
rect 5897 53830 5907 53882
rect 5931 53830 5961 53882
rect 5961 53830 5973 53882
rect 5973 53830 5987 53882
rect 6011 53830 6025 53882
rect 6025 53830 6037 53882
rect 6037 53830 6067 53882
rect 6091 53830 6101 53882
rect 6101 53830 6147 53882
rect 5851 53828 5907 53830
rect 5931 53828 5987 53830
rect 6011 53828 6067 53830
rect 6091 53828 6147 53830
rect 5851 52794 5907 52796
rect 5931 52794 5987 52796
rect 6011 52794 6067 52796
rect 6091 52794 6147 52796
rect 5851 52742 5897 52794
rect 5897 52742 5907 52794
rect 5931 52742 5961 52794
rect 5961 52742 5973 52794
rect 5973 52742 5987 52794
rect 6011 52742 6025 52794
rect 6025 52742 6037 52794
rect 6037 52742 6067 52794
rect 6091 52742 6101 52794
rect 6101 52742 6147 52794
rect 5851 52740 5907 52742
rect 5931 52740 5987 52742
rect 6011 52740 6067 52742
rect 6091 52740 6147 52742
rect 5851 51706 5907 51708
rect 5931 51706 5987 51708
rect 6011 51706 6067 51708
rect 6091 51706 6147 51708
rect 5851 51654 5897 51706
rect 5897 51654 5907 51706
rect 5931 51654 5961 51706
rect 5961 51654 5973 51706
rect 5973 51654 5987 51706
rect 6011 51654 6025 51706
rect 6025 51654 6037 51706
rect 6037 51654 6067 51706
rect 6091 51654 6101 51706
rect 6101 51654 6147 51706
rect 5851 51652 5907 51654
rect 5931 51652 5987 51654
rect 6011 51652 6067 51654
rect 6091 51652 6147 51654
rect 5814 51312 5870 51368
rect 5851 50618 5907 50620
rect 5931 50618 5987 50620
rect 6011 50618 6067 50620
rect 6091 50618 6147 50620
rect 5851 50566 5897 50618
rect 5897 50566 5907 50618
rect 5931 50566 5961 50618
rect 5961 50566 5973 50618
rect 5973 50566 5987 50618
rect 6011 50566 6025 50618
rect 6025 50566 6037 50618
rect 6037 50566 6067 50618
rect 6091 50566 6101 50618
rect 6101 50566 6147 50618
rect 5851 50564 5907 50566
rect 5931 50564 5987 50566
rect 6011 50564 6067 50566
rect 6091 50564 6147 50566
rect 5851 49530 5907 49532
rect 5931 49530 5987 49532
rect 6011 49530 6067 49532
rect 6091 49530 6147 49532
rect 5851 49478 5897 49530
rect 5897 49478 5907 49530
rect 5931 49478 5961 49530
rect 5961 49478 5973 49530
rect 5973 49478 5987 49530
rect 6011 49478 6025 49530
rect 6025 49478 6037 49530
rect 6037 49478 6067 49530
rect 6091 49478 6101 49530
rect 6101 49478 6147 49530
rect 5851 49476 5907 49478
rect 5931 49476 5987 49478
rect 6011 49476 6067 49478
rect 6091 49476 6147 49478
rect 5851 48442 5907 48444
rect 5931 48442 5987 48444
rect 6011 48442 6067 48444
rect 6091 48442 6147 48444
rect 5851 48390 5897 48442
rect 5897 48390 5907 48442
rect 5931 48390 5961 48442
rect 5961 48390 5973 48442
rect 5973 48390 5987 48442
rect 6011 48390 6025 48442
rect 6025 48390 6037 48442
rect 6037 48390 6067 48442
rect 6091 48390 6101 48442
rect 6101 48390 6147 48442
rect 5851 48388 5907 48390
rect 5931 48388 5987 48390
rect 6011 48388 6067 48390
rect 6091 48388 6147 48390
rect 5851 47354 5907 47356
rect 5931 47354 5987 47356
rect 6011 47354 6067 47356
rect 6091 47354 6147 47356
rect 5851 47302 5897 47354
rect 5897 47302 5907 47354
rect 5931 47302 5961 47354
rect 5961 47302 5973 47354
rect 5973 47302 5987 47354
rect 6011 47302 6025 47354
rect 6025 47302 6037 47354
rect 6037 47302 6067 47354
rect 6091 47302 6101 47354
rect 6101 47302 6147 47354
rect 5851 47300 5907 47302
rect 5931 47300 5987 47302
rect 6011 47300 6067 47302
rect 6091 47300 6147 47302
rect 5851 46266 5907 46268
rect 5931 46266 5987 46268
rect 6011 46266 6067 46268
rect 6091 46266 6147 46268
rect 5851 46214 5897 46266
rect 5897 46214 5907 46266
rect 5931 46214 5961 46266
rect 5961 46214 5973 46266
rect 5973 46214 5987 46266
rect 6011 46214 6025 46266
rect 6025 46214 6037 46266
rect 6037 46214 6067 46266
rect 6091 46214 6101 46266
rect 6101 46214 6147 46266
rect 5851 46212 5907 46214
rect 5931 46212 5987 46214
rect 6011 46212 6067 46214
rect 6091 46212 6147 46214
rect 5851 45178 5907 45180
rect 5931 45178 5987 45180
rect 6011 45178 6067 45180
rect 6091 45178 6147 45180
rect 5851 45126 5897 45178
rect 5897 45126 5907 45178
rect 5931 45126 5961 45178
rect 5961 45126 5973 45178
rect 5973 45126 5987 45178
rect 6011 45126 6025 45178
rect 6025 45126 6037 45178
rect 6037 45126 6067 45178
rect 6091 45126 6101 45178
rect 6101 45126 6147 45178
rect 5851 45124 5907 45126
rect 5931 45124 5987 45126
rect 6011 45124 6067 45126
rect 6091 45124 6147 45126
rect 5851 44090 5907 44092
rect 5931 44090 5987 44092
rect 6011 44090 6067 44092
rect 6091 44090 6147 44092
rect 5851 44038 5897 44090
rect 5897 44038 5907 44090
rect 5931 44038 5961 44090
rect 5961 44038 5973 44090
rect 5973 44038 5987 44090
rect 6011 44038 6025 44090
rect 6025 44038 6037 44090
rect 6037 44038 6067 44090
rect 6091 44038 6101 44090
rect 6101 44038 6147 44090
rect 5851 44036 5907 44038
rect 5931 44036 5987 44038
rect 6011 44036 6067 44038
rect 6091 44036 6147 44038
rect 5851 43002 5907 43004
rect 5931 43002 5987 43004
rect 6011 43002 6067 43004
rect 6091 43002 6147 43004
rect 5851 42950 5897 43002
rect 5897 42950 5907 43002
rect 5931 42950 5961 43002
rect 5961 42950 5973 43002
rect 5973 42950 5987 43002
rect 6011 42950 6025 43002
rect 6025 42950 6037 43002
rect 6037 42950 6067 43002
rect 6091 42950 6101 43002
rect 6101 42950 6147 43002
rect 5851 42948 5907 42950
rect 5931 42948 5987 42950
rect 6011 42948 6067 42950
rect 6091 42948 6147 42950
rect 5851 41914 5907 41916
rect 5931 41914 5987 41916
rect 6011 41914 6067 41916
rect 6091 41914 6147 41916
rect 5851 41862 5897 41914
rect 5897 41862 5907 41914
rect 5931 41862 5961 41914
rect 5961 41862 5973 41914
rect 5973 41862 5987 41914
rect 6011 41862 6025 41914
rect 6025 41862 6037 41914
rect 6037 41862 6067 41914
rect 6091 41862 6101 41914
rect 6101 41862 6147 41914
rect 5851 41860 5907 41862
rect 5931 41860 5987 41862
rect 6011 41860 6067 41862
rect 6091 41860 6147 41862
rect 5851 40826 5907 40828
rect 5931 40826 5987 40828
rect 6011 40826 6067 40828
rect 6091 40826 6147 40828
rect 5851 40774 5897 40826
rect 5897 40774 5907 40826
rect 5931 40774 5961 40826
rect 5961 40774 5973 40826
rect 5973 40774 5987 40826
rect 6011 40774 6025 40826
rect 6025 40774 6037 40826
rect 6037 40774 6067 40826
rect 6091 40774 6101 40826
rect 6101 40774 6147 40826
rect 5851 40772 5907 40774
rect 5931 40772 5987 40774
rect 6011 40772 6067 40774
rect 6091 40772 6147 40774
rect 5851 39738 5907 39740
rect 5931 39738 5987 39740
rect 6011 39738 6067 39740
rect 6091 39738 6147 39740
rect 5851 39686 5897 39738
rect 5897 39686 5907 39738
rect 5931 39686 5961 39738
rect 5961 39686 5973 39738
rect 5973 39686 5987 39738
rect 6011 39686 6025 39738
rect 6025 39686 6037 39738
rect 6037 39686 6067 39738
rect 6091 39686 6101 39738
rect 6101 39686 6147 39738
rect 5851 39684 5907 39686
rect 5931 39684 5987 39686
rect 6011 39684 6067 39686
rect 6091 39684 6147 39686
rect 5851 38650 5907 38652
rect 5931 38650 5987 38652
rect 6011 38650 6067 38652
rect 6091 38650 6147 38652
rect 5851 38598 5897 38650
rect 5897 38598 5907 38650
rect 5931 38598 5961 38650
rect 5961 38598 5973 38650
rect 5973 38598 5987 38650
rect 6011 38598 6025 38650
rect 6025 38598 6037 38650
rect 6037 38598 6067 38650
rect 6091 38598 6101 38650
rect 6101 38598 6147 38650
rect 5851 38596 5907 38598
rect 5931 38596 5987 38598
rect 6011 38596 6067 38598
rect 6091 38596 6147 38598
rect 5851 37562 5907 37564
rect 5931 37562 5987 37564
rect 6011 37562 6067 37564
rect 6091 37562 6147 37564
rect 5851 37510 5897 37562
rect 5897 37510 5907 37562
rect 5931 37510 5961 37562
rect 5961 37510 5973 37562
rect 5973 37510 5987 37562
rect 6011 37510 6025 37562
rect 6025 37510 6037 37562
rect 6037 37510 6067 37562
rect 6091 37510 6101 37562
rect 6101 37510 6147 37562
rect 5851 37508 5907 37510
rect 5931 37508 5987 37510
rect 6011 37508 6067 37510
rect 6091 37508 6147 37510
rect 5851 36474 5907 36476
rect 5931 36474 5987 36476
rect 6011 36474 6067 36476
rect 6091 36474 6147 36476
rect 5851 36422 5897 36474
rect 5897 36422 5907 36474
rect 5931 36422 5961 36474
rect 5961 36422 5973 36474
rect 5973 36422 5987 36474
rect 6011 36422 6025 36474
rect 6025 36422 6037 36474
rect 6037 36422 6067 36474
rect 6091 36422 6101 36474
rect 6101 36422 6147 36474
rect 5851 36420 5907 36422
rect 5931 36420 5987 36422
rect 6011 36420 6067 36422
rect 6091 36420 6147 36422
rect 5851 35386 5907 35388
rect 5931 35386 5987 35388
rect 6011 35386 6067 35388
rect 6091 35386 6147 35388
rect 5851 35334 5897 35386
rect 5897 35334 5907 35386
rect 5931 35334 5961 35386
rect 5961 35334 5973 35386
rect 5973 35334 5987 35386
rect 6011 35334 6025 35386
rect 6025 35334 6037 35386
rect 6037 35334 6067 35386
rect 6091 35334 6101 35386
rect 6101 35334 6147 35386
rect 5851 35332 5907 35334
rect 5931 35332 5987 35334
rect 6011 35332 6067 35334
rect 6091 35332 6147 35334
rect 5851 34298 5907 34300
rect 5931 34298 5987 34300
rect 6011 34298 6067 34300
rect 6091 34298 6147 34300
rect 5851 34246 5897 34298
rect 5897 34246 5907 34298
rect 5931 34246 5961 34298
rect 5961 34246 5973 34298
rect 5973 34246 5987 34298
rect 6011 34246 6025 34298
rect 6025 34246 6037 34298
rect 6037 34246 6067 34298
rect 6091 34246 6101 34298
rect 6101 34246 6147 34298
rect 5851 34244 5907 34246
rect 5931 34244 5987 34246
rect 6011 34244 6067 34246
rect 6091 34244 6147 34246
rect 5851 33210 5907 33212
rect 5931 33210 5987 33212
rect 6011 33210 6067 33212
rect 6091 33210 6147 33212
rect 5851 33158 5897 33210
rect 5897 33158 5907 33210
rect 5931 33158 5961 33210
rect 5961 33158 5973 33210
rect 5973 33158 5987 33210
rect 6011 33158 6025 33210
rect 6025 33158 6037 33210
rect 6037 33158 6067 33210
rect 6091 33158 6101 33210
rect 6101 33158 6147 33210
rect 5851 33156 5907 33158
rect 5931 33156 5987 33158
rect 6011 33156 6067 33158
rect 6091 33156 6147 33158
rect 5851 32122 5907 32124
rect 5931 32122 5987 32124
rect 6011 32122 6067 32124
rect 6091 32122 6147 32124
rect 5851 32070 5897 32122
rect 5897 32070 5907 32122
rect 5931 32070 5961 32122
rect 5961 32070 5973 32122
rect 5973 32070 5987 32122
rect 6011 32070 6025 32122
rect 6025 32070 6037 32122
rect 6037 32070 6067 32122
rect 6091 32070 6101 32122
rect 6101 32070 6147 32122
rect 5851 32068 5907 32070
rect 5931 32068 5987 32070
rect 6011 32068 6067 32070
rect 6091 32068 6147 32070
rect 5851 31034 5907 31036
rect 5931 31034 5987 31036
rect 6011 31034 6067 31036
rect 6091 31034 6147 31036
rect 5851 30982 5897 31034
rect 5897 30982 5907 31034
rect 5931 30982 5961 31034
rect 5961 30982 5973 31034
rect 5973 30982 5987 31034
rect 6011 30982 6025 31034
rect 6025 30982 6037 31034
rect 6037 30982 6067 31034
rect 6091 30982 6101 31034
rect 6101 30982 6147 31034
rect 5851 30980 5907 30982
rect 5931 30980 5987 30982
rect 6011 30980 6067 30982
rect 6091 30980 6147 30982
rect 5851 29946 5907 29948
rect 5931 29946 5987 29948
rect 6011 29946 6067 29948
rect 6091 29946 6147 29948
rect 5851 29894 5897 29946
rect 5897 29894 5907 29946
rect 5931 29894 5961 29946
rect 5961 29894 5973 29946
rect 5973 29894 5987 29946
rect 6011 29894 6025 29946
rect 6025 29894 6037 29946
rect 6037 29894 6067 29946
rect 6091 29894 6101 29946
rect 6101 29894 6147 29946
rect 5851 29892 5907 29894
rect 5931 29892 5987 29894
rect 6011 29892 6067 29894
rect 6091 29892 6147 29894
rect 5851 28858 5907 28860
rect 5931 28858 5987 28860
rect 6011 28858 6067 28860
rect 6091 28858 6147 28860
rect 5851 28806 5897 28858
rect 5897 28806 5907 28858
rect 5931 28806 5961 28858
rect 5961 28806 5973 28858
rect 5973 28806 5987 28858
rect 6011 28806 6025 28858
rect 6025 28806 6037 28858
rect 6037 28806 6067 28858
rect 6091 28806 6101 28858
rect 6101 28806 6147 28858
rect 5851 28804 5907 28806
rect 5931 28804 5987 28806
rect 6011 28804 6067 28806
rect 6091 28804 6147 28806
rect 5851 27770 5907 27772
rect 5931 27770 5987 27772
rect 6011 27770 6067 27772
rect 6091 27770 6147 27772
rect 5851 27718 5897 27770
rect 5897 27718 5907 27770
rect 5931 27718 5961 27770
rect 5961 27718 5973 27770
rect 5973 27718 5987 27770
rect 6011 27718 6025 27770
rect 6025 27718 6037 27770
rect 6037 27718 6067 27770
rect 6091 27718 6101 27770
rect 6101 27718 6147 27770
rect 5851 27716 5907 27718
rect 5931 27716 5987 27718
rect 6011 27716 6067 27718
rect 6091 27716 6147 27718
rect 5851 26682 5907 26684
rect 5931 26682 5987 26684
rect 6011 26682 6067 26684
rect 6091 26682 6147 26684
rect 5851 26630 5897 26682
rect 5897 26630 5907 26682
rect 5931 26630 5961 26682
rect 5961 26630 5973 26682
rect 5973 26630 5987 26682
rect 6011 26630 6025 26682
rect 6025 26630 6037 26682
rect 6037 26630 6067 26682
rect 6091 26630 6101 26682
rect 6101 26630 6147 26682
rect 5851 26628 5907 26630
rect 5931 26628 5987 26630
rect 6011 26628 6067 26630
rect 6091 26628 6147 26630
rect 5851 25594 5907 25596
rect 5931 25594 5987 25596
rect 6011 25594 6067 25596
rect 6091 25594 6147 25596
rect 5851 25542 5897 25594
rect 5897 25542 5907 25594
rect 5931 25542 5961 25594
rect 5961 25542 5973 25594
rect 5973 25542 5987 25594
rect 6011 25542 6025 25594
rect 6025 25542 6037 25594
rect 6037 25542 6067 25594
rect 6091 25542 6101 25594
rect 6101 25542 6147 25594
rect 5851 25540 5907 25542
rect 5931 25540 5987 25542
rect 6011 25540 6067 25542
rect 6091 25540 6147 25542
rect 5851 24506 5907 24508
rect 5931 24506 5987 24508
rect 6011 24506 6067 24508
rect 6091 24506 6147 24508
rect 5851 24454 5897 24506
rect 5897 24454 5907 24506
rect 5931 24454 5961 24506
rect 5961 24454 5973 24506
rect 5973 24454 5987 24506
rect 6011 24454 6025 24506
rect 6025 24454 6037 24506
rect 6037 24454 6067 24506
rect 6091 24454 6101 24506
rect 6101 24454 6147 24506
rect 5851 24452 5907 24454
rect 5931 24452 5987 24454
rect 6011 24452 6067 24454
rect 6091 24452 6147 24454
rect 5851 23418 5907 23420
rect 5931 23418 5987 23420
rect 6011 23418 6067 23420
rect 6091 23418 6147 23420
rect 5851 23366 5897 23418
rect 5897 23366 5907 23418
rect 5931 23366 5961 23418
rect 5961 23366 5973 23418
rect 5973 23366 5987 23418
rect 6011 23366 6025 23418
rect 6025 23366 6037 23418
rect 6037 23366 6067 23418
rect 6091 23366 6101 23418
rect 6101 23366 6147 23418
rect 5851 23364 5907 23366
rect 5931 23364 5987 23366
rect 6011 23364 6067 23366
rect 6091 23364 6147 23366
rect 5851 22330 5907 22332
rect 5931 22330 5987 22332
rect 6011 22330 6067 22332
rect 6091 22330 6147 22332
rect 5851 22278 5897 22330
rect 5897 22278 5907 22330
rect 5931 22278 5961 22330
rect 5961 22278 5973 22330
rect 5973 22278 5987 22330
rect 6011 22278 6025 22330
rect 6025 22278 6037 22330
rect 6037 22278 6067 22330
rect 6091 22278 6101 22330
rect 6101 22278 6147 22330
rect 5851 22276 5907 22278
rect 5931 22276 5987 22278
rect 6011 22276 6067 22278
rect 6091 22276 6147 22278
rect 5851 21242 5907 21244
rect 5931 21242 5987 21244
rect 6011 21242 6067 21244
rect 6091 21242 6147 21244
rect 5851 21190 5897 21242
rect 5897 21190 5907 21242
rect 5931 21190 5961 21242
rect 5961 21190 5973 21242
rect 5973 21190 5987 21242
rect 6011 21190 6025 21242
rect 6025 21190 6037 21242
rect 6037 21190 6067 21242
rect 6091 21190 6101 21242
rect 6101 21190 6147 21242
rect 5851 21188 5907 21190
rect 5931 21188 5987 21190
rect 6011 21188 6067 21190
rect 6091 21188 6147 21190
rect 5851 20154 5907 20156
rect 5931 20154 5987 20156
rect 6011 20154 6067 20156
rect 6091 20154 6147 20156
rect 5851 20102 5897 20154
rect 5897 20102 5907 20154
rect 5931 20102 5961 20154
rect 5961 20102 5973 20154
rect 5973 20102 5987 20154
rect 6011 20102 6025 20154
rect 6025 20102 6037 20154
rect 6037 20102 6067 20154
rect 6091 20102 6101 20154
rect 6101 20102 6147 20154
rect 5851 20100 5907 20102
rect 5931 20100 5987 20102
rect 6011 20100 6067 20102
rect 6091 20100 6147 20102
rect 5851 19066 5907 19068
rect 5931 19066 5987 19068
rect 6011 19066 6067 19068
rect 6091 19066 6147 19068
rect 5851 19014 5897 19066
rect 5897 19014 5907 19066
rect 5931 19014 5961 19066
rect 5961 19014 5973 19066
rect 5973 19014 5987 19066
rect 6011 19014 6025 19066
rect 6025 19014 6037 19066
rect 6037 19014 6067 19066
rect 6091 19014 6101 19066
rect 6101 19014 6147 19066
rect 5851 19012 5907 19014
rect 5931 19012 5987 19014
rect 6011 19012 6067 19014
rect 6091 19012 6147 19014
rect 5851 17978 5907 17980
rect 5931 17978 5987 17980
rect 6011 17978 6067 17980
rect 6091 17978 6147 17980
rect 5851 17926 5897 17978
rect 5897 17926 5907 17978
rect 5931 17926 5961 17978
rect 5961 17926 5973 17978
rect 5973 17926 5987 17978
rect 6011 17926 6025 17978
rect 6025 17926 6037 17978
rect 6037 17926 6067 17978
rect 6091 17926 6101 17978
rect 6101 17926 6147 17978
rect 5851 17924 5907 17926
rect 5931 17924 5987 17926
rect 6011 17924 6067 17926
rect 6091 17924 6147 17926
rect 5851 16890 5907 16892
rect 5931 16890 5987 16892
rect 6011 16890 6067 16892
rect 6091 16890 6147 16892
rect 5851 16838 5897 16890
rect 5897 16838 5907 16890
rect 5931 16838 5961 16890
rect 5961 16838 5973 16890
rect 5973 16838 5987 16890
rect 6011 16838 6025 16890
rect 6025 16838 6037 16890
rect 6037 16838 6067 16890
rect 6091 16838 6101 16890
rect 6101 16838 6147 16890
rect 5851 16836 5907 16838
rect 5931 16836 5987 16838
rect 6011 16836 6067 16838
rect 6091 16836 6147 16838
rect 5851 15802 5907 15804
rect 5931 15802 5987 15804
rect 6011 15802 6067 15804
rect 6091 15802 6147 15804
rect 5851 15750 5897 15802
rect 5897 15750 5907 15802
rect 5931 15750 5961 15802
rect 5961 15750 5973 15802
rect 5973 15750 5987 15802
rect 6011 15750 6025 15802
rect 6025 15750 6037 15802
rect 6037 15750 6067 15802
rect 6091 15750 6101 15802
rect 6101 15750 6147 15802
rect 5851 15748 5907 15750
rect 5931 15748 5987 15750
rect 6011 15748 6067 15750
rect 6091 15748 6147 15750
rect 7483 74010 7539 74012
rect 7563 74010 7619 74012
rect 7643 74010 7699 74012
rect 7723 74010 7779 74012
rect 7483 73958 7529 74010
rect 7529 73958 7539 74010
rect 7563 73958 7593 74010
rect 7593 73958 7605 74010
rect 7605 73958 7619 74010
rect 7643 73958 7657 74010
rect 7657 73958 7669 74010
rect 7669 73958 7699 74010
rect 7723 73958 7733 74010
rect 7733 73958 7779 74010
rect 7483 73956 7539 73958
rect 7563 73956 7619 73958
rect 7643 73956 7699 73958
rect 7723 73956 7779 73958
rect 9115 76730 9171 76732
rect 9195 76730 9251 76732
rect 9275 76730 9331 76732
rect 9355 76730 9411 76732
rect 9115 76678 9161 76730
rect 9161 76678 9171 76730
rect 9195 76678 9225 76730
rect 9225 76678 9237 76730
rect 9237 76678 9251 76730
rect 9275 76678 9289 76730
rect 9289 76678 9301 76730
rect 9301 76678 9331 76730
rect 9355 76678 9365 76730
rect 9365 76678 9411 76730
rect 9115 76676 9171 76678
rect 9195 76676 9251 76678
rect 9275 76676 9331 76678
rect 9355 76676 9411 76678
rect 9115 75642 9171 75644
rect 9195 75642 9251 75644
rect 9275 75642 9331 75644
rect 9355 75642 9411 75644
rect 9115 75590 9161 75642
rect 9161 75590 9171 75642
rect 9195 75590 9225 75642
rect 9225 75590 9237 75642
rect 9237 75590 9251 75642
rect 9275 75590 9289 75642
rect 9289 75590 9301 75642
rect 9301 75590 9331 75642
rect 9355 75590 9365 75642
rect 9365 75590 9411 75642
rect 9115 75588 9171 75590
rect 9195 75588 9251 75590
rect 9275 75588 9331 75590
rect 9355 75588 9411 75590
rect 9115 74554 9171 74556
rect 9195 74554 9251 74556
rect 9275 74554 9331 74556
rect 9355 74554 9411 74556
rect 9115 74502 9161 74554
rect 9161 74502 9171 74554
rect 9195 74502 9225 74554
rect 9225 74502 9237 74554
rect 9237 74502 9251 74554
rect 9275 74502 9289 74554
rect 9289 74502 9301 74554
rect 9301 74502 9331 74554
rect 9355 74502 9365 74554
rect 9365 74502 9411 74554
rect 9115 74500 9171 74502
rect 9195 74500 9251 74502
rect 9275 74500 9331 74502
rect 9355 74500 9411 74502
rect 10046 76472 10102 76528
rect 10046 75692 10048 75712
rect 10048 75692 10100 75712
rect 10100 75692 10102 75712
rect 10046 75656 10102 75692
rect 10046 74976 10102 75032
rect 10046 74160 10102 74216
rect 10046 73516 10048 73536
rect 10048 73516 10100 73536
rect 10100 73516 10102 73536
rect 10046 73480 10102 73516
rect 9115 73466 9171 73468
rect 9195 73466 9251 73468
rect 9275 73466 9331 73468
rect 9355 73466 9411 73468
rect 9115 73414 9161 73466
rect 9161 73414 9171 73466
rect 9195 73414 9225 73466
rect 9225 73414 9237 73466
rect 9237 73414 9251 73466
rect 9275 73414 9289 73466
rect 9289 73414 9301 73466
rect 9301 73414 9331 73466
rect 9355 73414 9365 73466
rect 9365 73414 9411 73466
rect 9115 73412 9171 73414
rect 9195 73412 9251 73414
rect 9275 73412 9331 73414
rect 9355 73412 9411 73414
rect 7483 72922 7539 72924
rect 7563 72922 7619 72924
rect 7643 72922 7699 72924
rect 7723 72922 7779 72924
rect 7483 72870 7529 72922
rect 7529 72870 7539 72922
rect 7563 72870 7593 72922
rect 7593 72870 7605 72922
rect 7605 72870 7619 72922
rect 7643 72870 7657 72922
rect 7657 72870 7669 72922
rect 7669 72870 7699 72922
rect 7723 72870 7733 72922
rect 7733 72870 7779 72922
rect 7483 72868 7539 72870
rect 7563 72868 7619 72870
rect 7643 72868 7699 72870
rect 7723 72868 7779 72870
rect 10046 72664 10102 72720
rect 6642 41248 6698 41304
rect 6458 36896 6514 36952
rect 9115 72378 9171 72380
rect 9195 72378 9251 72380
rect 9275 72378 9331 72380
rect 9355 72378 9411 72380
rect 9115 72326 9161 72378
rect 9161 72326 9171 72378
rect 9195 72326 9225 72378
rect 9225 72326 9237 72378
rect 9237 72326 9251 72378
rect 9275 72326 9289 72378
rect 9289 72326 9301 72378
rect 9301 72326 9331 72378
rect 9355 72326 9365 72378
rect 9365 72326 9411 72378
rect 9115 72324 9171 72326
rect 9195 72324 9251 72326
rect 9275 72324 9331 72326
rect 9355 72324 9411 72326
rect 10046 71884 10048 71904
rect 10048 71884 10100 71904
rect 10100 71884 10102 71904
rect 7483 71834 7539 71836
rect 7563 71834 7619 71836
rect 7643 71834 7699 71836
rect 7723 71834 7779 71836
rect 7483 71782 7529 71834
rect 7529 71782 7539 71834
rect 7563 71782 7593 71834
rect 7593 71782 7605 71834
rect 7605 71782 7619 71834
rect 7643 71782 7657 71834
rect 7657 71782 7669 71834
rect 7669 71782 7699 71834
rect 7723 71782 7733 71834
rect 7733 71782 7779 71834
rect 7483 71780 7539 71782
rect 7563 71780 7619 71782
rect 7643 71780 7699 71782
rect 7723 71780 7779 71782
rect 10046 71848 10102 71884
rect 9115 71290 9171 71292
rect 9195 71290 9251 71292
rect 9275 71290 9331 71292
rect 9355 71290 9411 71292
rect 9115 71238 9161 71290
rect 9161 71238 9171 71290
rect 9195 71238 9225 71290
rect 9225 71238 9237 71290
rect 9237 71238 9251 71290
rect 9275 71238 9289 71290
rect 9289 71238 9301 71290
rect 9301 71238 9331 71290
rect 9355 71238 9365 71290
rect 9365 71238 9411 71290
rect 9115 71236 9171 71238
rect 9195 71236 9251 71238
rect 9275 71236 9331 71238
rect 9355 71236 9411 71238
rect 7483 70746 7539 70748
rect 7563 70746 7619 70748
rect 7643 70746 7699 70748
rect 7723 70746 7779 70748
rect 7483 70694 7529 70746
rect 7529 70694 7539 70746
rect 7563 70694 7593 70746
rect 7593 70694 7605 70746
rect 7605 70694 7619 70746
rect 7643 70694 7657 70746
rect 7657 70694 7669 70746
rect 7669 70694 7699 70746
rect 7723 70694 7733 70746
rect 7733 70694 7779 70746
rect 7483 70692 7539 70694
rect 7563 70692 7619 70694
rect 7643 70692 7699 70694
rect 7723 70692 7779 70694
rect 10046 71168 10102 71224
rect 10690 70352 10746 70408
rect 9115 70202 9171 70204
rect 9195 70202 9251 70204
rect 9275 70202 9331 70204
rect 9355 70202 9411 70204
rect 9115 70150 9161 70202
rect 9161 70150 9171 70202
rect 9195 70150 9225 70202
rect 9225 70150 9237 70202
rect 9237 70150 9251 70202
rect 9275 70150 9289 70202
rect 9289 70150 9301 70202
rect 9301 70150 9331 70202
rect 9355 70150 9365 70202
rect 9365 70150 9411 70202
rect 9115 70148 9171 70150
rect 9195 70148 9251 70150
rect 9275 70148 9331 70150
rect 9355 70148 9411 70150
rect 10046 69708 10048 69728
rect 10048 69708 10100 69728
rect 10100 69708 10102 69728
rect 10046 69672 10102 69708
rect 7483 69658 7539 69660
rect 7563 69658 7619 69660
rect 7643 69658 7699 69660
rect 7723 69658 7779 69660
rect 7483 69606 7529 69658
rect 7529 69606 7539 69658
rect 7563 69606 7593 69658
rect 7593 69606 7605 69658
rect 7605 69606 7619 69658
rect 7643 69606 7657 69658
rect 7657 69606 7669 69658
rect 7669 69606 7699 69658
rect 7723 69606 7733 69658
rect 7733 69606 7779 69658
rect 7483 69604 7539 69606
rect 7563 69604 7619 69606
rect 7643 69604 7699 69606
rect 7723 69604 7779 69606
rect 9115 69114 9171 69116
rect 9195 69114 9251 69116
rect 9275 69114 9331 69116
rect 9355 69114 9411 69116
rect 9115 69062 9161 69114
rect 9161 69062 9171 69114
rect 9195 69062 9225 69114
rect 9225 69062 9237 69114
rect 9237 69062 9251 69114
rect 9275 69062 9289 69114
rect 9289 69062 9301 69114
rect 9301 69062 9331 69114
rect 9355 69062 9365 69114
rect 9365 69062 9411 69114
rect 9115 69060 9171 69062
rect 9195 69060 9251 69062
rect 9275 69060 9331 69062
rect 9355 69060 9411 69062
rect 10046 68856 10102 68912
rect 7483 68570 7539 68572
rect 7563 68570 7619 68572
rect 7643 68570 7699 68572
rect 7723 68570 7779 68572
rect 7483 68518 7529 68570
rect 7529 68518 7539 68570
rect 7563 68518 7593 68570
rect 7593 68518 7605 68570
rect 7605 68518 7619 68570
rect 7643 68518 7657 68570
rect 7657 68518 7669 68570
rect 7669 68518 7699 68570
rect 7723 68518 7733 68570
rect 7733 68518 7779 68570
rect 7483 68516 7539 68518
rect 7563 68516 7619 68518
rect 7643 68516 7699 68518
rect 7723 68516 7779 68518
rect 9115 68026 9171 68028
rect 9195 68026 9251 68028
rect 9275 68026 9331 68028
rect 9355 68026 9411 68028
rect 9115 67974 9161 68026
rect 9161 67974 9171 68026
rect 9195 67974 9225 68026
rect 9225 67974 9237 68026
rect 9237 67974 9251 68026
rect 9275 67974 9289 68026
rect 9289 67974 9301 68026
rect 9301 67974 9331 68026
rect 9355 67974 9365 68026
rect 9365 67974 9411 68026
rect 9115 67972 9171 67974
rect 9195 67972 9251 67974
rect 9275 67972 9331 67974
rect 9355 67972 9411 67974
rect 7483 67482 7539 67484
rect 7563 67482 7619 67484
rect 7643 67482 7699 67484
rect 7723 67482 7779 67484
rect 7483 67430 7529 67482
rect 7529 67430 7539 67482
rect 7563 67430 7593 67482
rect 7593 67430 7605 67482
rect 7605 67430 7619 67482
rect 7643 67430 7657 67482
rect 7657 67430 7669 67482
rect 7669 67430 7699 67482
rect 7723 67430 7733 67482
rect 7733 67430 7779 67482
rect 7483 67428 7539 67430
rect 7563 67428 7619 67430
rect 7643 67428 7699 67430
rect 7723 67428 7779 67430
rect 9115 66938 9171 66940
rect 9195 66938 9251 66940
rect 9275 66938 9331 66940
rect 9355 66938 9411 66940
rect 9115 66886 9161 66938
rect 9161 66886 9171 66938
rect 9195 66886 9225 66938
rect 9225 66886 9237 66938
rect 9237 66886 9251 66938
rect 9275 66886 9289 66938
rect 9289 66886 9301 66938
rect 9301 66886 9331 66938
rect 9355 66886 9365 66938
rect 9365 66886 9411 66938
rect 9115 66884 9171 66886
rect 9195 66884 9251 66886
rect 9275 66884 9331 66886
rect 9355 66884 9411 66886
rect 7483 66394 7539 66396
rect 7563 66394 7619 66396
rect 7643 66394 7699 66396
rect 7723 66394 7779 66396
rect 7483 66342 7529 66394
rect 7529 66342 7539 66394
rect 7563 66342 7593 66394
rect 7593 66342 7605 66394
rect 7605 66342 7619 66394
rect 7643 66342 7657 66394
rect 7657 66342 7669 66394
rect 7669 66342 7699 66394
rect 7723 66342 7733 66394
rect 7733 66342 7779 66394
rect 7483 66340 7539 66342
rect 7563 66340 7619 66342
rect 7643 66340 7699 66342
rect 7723 66340 7779 66342
rect 9115 65850 9171 65852
rect 9195 65850 9251 65852
rect 9275 65850 9331 65852
rect 9355 65850 9411 65852
rect 9115 65798 9161 65850
rect 9161 65798 9171 65850
rect 9195 65798 9225 65850
rect 9225 65798 9237 65850
rect 9237 65798 9251 65850
rect 9275 65798 9289 65850
rect 9289 65798 9301 65850
rect 9301 65798 9331 65850
rect 9355 65798 9365 65850
rect 9365 65798 9411 65850
rect 9115 65796 9171 65798
rect 9195 65796 9251 65798
rect 9275 65796 9331 65798
rect 9355 65796 9411 65798
rect 7483 65306 7539 65308
rect 7563 65306 7619 65308
rect 7643 65306 7699 65308
rect 7723 65306 7779 65308
rect 7483 65254 7529 65306
rect 7529 65254 7539 65306
rect 7563 65254 7593 65306
rect 7593 65254 7605 65306
rect 7605 65254 7619 65306
rect 7643 65254 7657 65306
rect 7657 65254 7669 65306
rect 7669 65254 7699 65306
rect 7723 65254 7733 65306
rect 7733 65254 7779 65306
rect 7483 65252 7539 65254
rect 7563 65252 7619 65254
rect 7643 65252 7699 65254
rect 7723 65252 7779 65254
rect 9115 64762 9171 64764
rect 9195 64762 9251 64764
rect 9275 64762 9331 64764
rect 9355 64762 9411 64764
rect 9115 64710 9161 64762
rect 9161 64710 9171 64762
rect 9195 64710 9225 64762
rect 9225 64710 9237 64762
rect 9237 64710 9251 64762
rect 9275 64710 9289 64762
rect 9289 64710 9301 64762
rect 9301 64710 9331 64762
rect 9355 64710 9365 64762
rect 9365 64710 9411 64762
rect 9115 64708 9171 64710
rect 9195 64708 9251 64710
rect 9275 64708 9331 64710
rect 9355 64708 9411 64710
rect 7483 64218 7539 64220
rect 7563 64218 7619 64220
rect 7643 64218 7699 64220
rect 7723 64218 7779 64220
rect 7483 64166 7529 64218
rect 7529 64166 7539 64218
rect 7563 64166 7593 64218
rect 7593 64166 7605 64218
rect 7605 64166 7619 64218
rect 7643 64166 7657 64218
rect 7657 64166 7669 64218
rect 7669 64166 7699 64218
rect 7723 64166 7733 64218
rect 7733 64166 7779 64218
rect 7483 64164 7539 64166
rect 7563 64164 7619 64166
rect 7643 64164 7699 64166
rect 7723 64164 7779 64166
rect 10046 68196 10102 68232
rect 10046 68176 10048 68196
rect 10048 68176 10100 68196
rect 10100 68176 10102 68196
rect 10046 67360 10102 67416
rect 10046 66680 10102 66736
rect 10046 65900 10048 65920
rect 10048 65900 10100 65920
rect 10100 65900 10102 65920
rect 10046 65864 10102 65900
rect 10046 65184 10102 65240
rect 7483 63130 7539 63132
rect 7563 63130 7619 63132
rect 7643 63130 7699 63132
rect 7723 63130 7779 63132
rect 7483 63078 7529 63130
rect 7529 63078 7539 63130
rect 7563 63078 7593 63130
rect 7593 63078 7605 63130
rect 7605 63078 7619 63130
rect 7643 63078 7657 63130
rect 7657 63078 7669 63130
rect 7669 63078 7699 63130
rect 7723 63078 7733 63130
rect 7733 63078 7779 63130
rect 7483 63076 7539 63078
rect 7563 63076 7619 63078
rect 7643 63076 7699 63078
rect 7723 63076 7779 63078
rect 7483 62042 7539 62044
rect 7563 62042 7619 62044
rect 7643 62042 7699 62044
rect 7723 62042 7779 62044
rect 7483 61990 7529 62042
rect 7529 61990 7539 62042
rect 7563 61990 7593 62042
rect 7593 61990 7605 62042
rect 7605 61990 7619 62042
rect 7643 61990 7657 62042
rect 7657 61990 7669 62042
rect 7669 61990 7699 62042
rect 7723 61990 7733 62042
rect 7733 61990 7779 62042
rect 7483 61988 7539 61990
rect 7563 61988 7619 61990
rect 7643 61988 7699 61990
rect 7723 61988 7779 61990
rect 7483 60954 7539 60956
rect 7563 60954 7619 60956
rect 7643 60954 7699 60956
rect 7723 60954 7779 60956
rect 7483 60902 7529 60954
rect 7529 60902 7539 60954
rect 7563 60902 7593 60954
rect 7593 60902 7605 60954
rect 7605 60902 7619 60954
rect 7643 60902 7657 60954
rect 7657 60902 7669 60954
rect 7669 60902 7699 60954
rect 7723 60902 7733 60954
rect 7733 60902 7779 60954
rect 7483 60900 7539 60902
rect 7563 60900 7619 60902
rect 7643 60900 7699 60902
rect 7723 60900 7779 60902
rect 7483 59866 7539 59868
rect 7563 59866 7619 59868
rect 7643 59866 7699 59868
rect 7723 59866 7779 59868
rect 7483 59814 7529 59866
rect 7529 59814 7539 59866
rect 7563 59814 7593 59866
rect 7593 59814 7605 59866
rect 7605 59814 7619 59866
rect 7643 59814 7657 59866
rect 7657 59814 7669 59866
rect 7669 59814 7699 59866
rect 7723 59814 7733 59866
rect 7733 59814 7779 59866
rect 7483 59812 7539 59814
rect 7563 59812 7619 59814
rect 7643 59812 7699 59814
rect 7723 59812 7779 59814
rect 7483 58778 7539 58780
rect 7563 58778 7619 58780
rect 7643 58778 7699 58780
rect 7723 58778 7779 58780
rect 7483 58726 7529 58778
rect 7529 58726 7539 58778
rect 7563 58726 7593 58778
rect 7593 58726 7605 58778
rect 7605 58726 7619 58778
rect 7643 58726 7657 58778
rect 7657 58726 7669 58778
rect 7669 58726 7699 58778
rect 7723 58726 7733 58778
rect 7733 58726 7779 58778
rect 7483 58724 7539 58726
rect 7563 58724 7619 58726
rect 7643 58724 7699 58726
rect 7723 58724 7779 58726
rect 7483 57690 7539 57692
rect 7563 57690 7619 57692
rect 7643 57690 7699 57692
rect 7723 57690 7779 57692
rect 7483 57638 7529 57690
rect 7529 57638 7539 57690
rect 7563 57638 7593 57690
rect 7593 57638 7605 57690
rect 7605 57638 7619 57690
rect 7643 57638 7657 57690
rect 7657 57638 7669 57690
rect 7669 57638 7699 57690
rect 7723 57638 7733 57690
rect 7733 57638 7779 57690
rect 7483 57636 7539 57638
rect 7563 57636 7619 57638
rect 7643 57636 7699 57638
rect 7723 57636 7779 57638
rect 7483 56602 7539 56604
rect 7563 56602 7619 56604
rect 7643 56602 7699 56604
rect 7723 56602 7779 56604
rect 7483 56550 7529 56602
rect 7529 56550 7539 56602
rect 7563 56550 7593 56602
rect 7593 56550 7605 56602
rect 7605 56550 7619 56602
rect 7643 56550 7657 56602
rect 7657 56550 7669 56602
rect 7669 56550 7699 56602
rect 7723 56550 7733 56602
rect 7733 56550 7779 56602
rect 7483 56548 7539 56550
rect 7563 56548 7619 56550
rect 7643 56548 7699 56550
rect 7723 56548 7779 56550
rect 7483 55514 7539 55516
rect 7563 55514 7619 55516
rect 7643 55514 7699 55516
rect 7723 55514 7779 55516
rect 7483 55462 7529 55514
rect 7529 55462 7539 55514
rect 7563 55462 7593 55514
rect 7593 55462 7605 55514
rect 7605 55462 7619 55514
rect 7643 55462 7657 55514
rect 7657 55462 7669 55514
rect 7669 55462 7699 55514
rect 7723 55462 7733 55514
rect 7733 55462 7779 55514
rect 7483 55460 7539 55462
rect 7563 55460 7619 55462
rect 7643 55460 7699 55462
rect 7723 55460 7779 55462
rect 7483 54426 7539 54428
rect 7563 54426 7619 54428
rect 7643 54426 7699 54428
rect 7723 54426 7779 54428
rect 7483 54374 7529 54426
rect 7529 54374 7539 54426
rect 7563 54374 7593 54426
rect 7593 54374 7605 54426
rect 7605 54374 7619 54426
rect 7643 54374 7657 54426
rect 7657 54374 7669 54426
rect 7669 54374 7699 54426
rect 7723 54374 7733 54426
rect 7733 54374 7779 54426
rect 7483 54372 7539 54374
rect 7563 54372 7619 54374
rect 7643 54372 7699 54374
rect 7723 54372 7779 54374
rect 7483 53338 7539 53340
rect 7563 53338 7619 53340
rect 7643 53338 7699 53340
rect 7723 53338 7779 53340
rect 7483 53286 7529 53338
rect 7529 53286 7539 53338
rect 7563 53286 7593 53338
rect 7593 53286 7605 53338
rect 7605 53286 7619 53338
rect 7643 53286 7657 53338
rect 7657 53286 7669 53338
rect 7669 53286 7699 53338
rect 7723 53286 7733 53338
rect 7733 53286 7779 53338
rect 7483 53284 7539 53286
rect 7563 53284 7619 53286
rect 7643 53284 7699 53286
rect 7723 53284 7779 53286
rect 7483 52250 7539 52252
rect 7563 52250 7619 52252
rect 7643 52250 7699 52252
rect 7723 52250 7779 52252
rect 7483 52198 7529 52250
rect 7529 52198 7539 52250
rect 7563 52198 7593 52250
rect 7593 52198 7605 52250
rect 7605 52198 7619 52250
rect 7643 52198 7657 52250
rect 7657 52198 7669 52250
rect 7669 52198 7699 52250
rect 7723 52198 7733 52250
rect 7733 52198 7779 52250
rect 7483 52196 7539 52198
rect 7563 52196 7619 52198
rect 7643 52196 7699 52198
rect 7723 52196 7779 52198
rect 7838 51448 7894 51504
rect 7483 51162 7539 51164
rect 7563 51162 7619 51164
rect 7643 51162 7699 51164
rect 7723 51162 7779 51164
rect 7483 51110 7529 51162
rect 7529 51110 7539 51162
rect 7563 51110 7593 51162
rect 7593 51110 7605 51162
rect 7605 51110 7619 51162
rect 7643 51110 7657 51162
rect 7657 51110 7669 51162
rect 7669 51110 7699 51162
rect 7723 51110 7733 51162
rect 7733 51110 7779 51162
rect 7483 51108 7539 51110
rect 7563 51108 7619 51110
rect 7643 51108 7699 51110
rect 7723 51108 7779 51110
rect 7483 50074 7539 50076
rect 7563 50074 7619 50076
rect 7643 50074 7699 50076
rect 7723 50074 7779 50076
rect 7483 50022 7529 50074
rect 7529 50022 7539 50074
rect 7563 50022 7593 50074
rect 7593 50022 7605 50074
rect 7605 50022 7619 50074
rect 7643 50022 7657 50074
rect 7657 50022 7669 50074
rect 7669 50022 7699 50074
rect 7723 50022 7733 50074
rect 7733 50022 7779 50074
rect 7483 50020 7539 50022
rect 7563 50020 7619 50022
rect 7643 50020 7699 50022
rect 7723 50020 7779 50022
rect 7483 48986 7539 48988
rect 7563 48986 7619 48988
rect 7643 48986 7699 48988
rect 7723 48986 7779 48988
rect 7483 48934 7529 48986
rect 7529 48934 7539 48986
rect 7563 48934 7593 48986
rect 7593 48934 7605 48986
rect 7605 48934 7619 48986
rect 7643 48934 7657 48986
rect 7657 48934 7669 48986
rect 7669 48934 7699 48986
rect 7723 48934 7733 48986
rect 7733 48934 7779 48986
rect 7483 48932 7539 48934
rect 7563 48932 7619 48934
rect 7643 48932 7699 48934
rect 7723 48932 7779 48934
rect 7483 47898 7539 47900
rect 7563 47898 7619 47900
rect 7643 47898 7699 47900
rect 7723 47898 7779 47900
rect 7483 47846 7529 47898
rect 7529 47846 7539 47898
rect 7563 47846 7593 47898
rect 7593 47846 7605 47898
rect 7605 47846 7619 47898
rect 7643 47846 7657 47898
rect 7657 47846 7669 47898
rect 7669 47846 7699 47898
rect 7723 47846 7733 47898
rect 7733 47846 7779 47898
rect 7483 47844 7539 47846
rect 7563 47844 7619 47846
rect 7643 47844 7699 47846
rect 7723 47844 7779 47846
rect 7483 46810 7539 46812
rect 7563 46810 7619 46812
rect 7643 46810 7699 46812
rect 7723 46810 7779 46812
rect 7483 46758 7529 46810
rect 7529 46758 7539 46810
rect 7563 46758 7593 46810
rect 7593 46758 7605 46810
rect 7605 46758 7619 46810
rect 7643 46758 7657 46810
rect 7657 46758 7669 46810
rect 7669 46758 7699 46810
rect 7723 46758 7733 46810
rect 7733 46758 7779 46810
rect 7483 46756 7539 46758
rect 7563 46756 7619 46758
rect 7643 46756 7699 46758
rect 7723 46756 7779 46758
rect 7483 45722 7539 45724
rect 7563 45722 7619 45724
rect 7643 45722 7699 45724
rect 7723 45722 7779 45724
rect 7483 45670 7529 45722
rect 7529 45670 7539 45722
rect 7563 45670 7593 45722
rect 7593 45670 7605 45722
rect 7605 45670 7619 45722
rect 7643 45670 7657 45722
rect 7657 45670 7669 45722
rect 7669 45670 7699 45722
rect 7723 45670 7733 45722
rect 7733 45670 7779 45722
rect 7483 45668 7539 45670
rect 7563 45668 7619 45670
rect 7643 45668 7699 45670
rect 7723 45668 7779 45670
rect 7483 44634 7539 44636
rect 7563 44634 7619 44636
rect 7643 44634 7699 44636
rect 7723 44634 7779 44636
rect 7483 44582 7529 44634
rect 7529 44582 7539 44634
rect 7563 44582 7593 44634
rect 7593 44582 7605 44634
rect 7605 44582 7619 44634
rect 7643 44582 7657 44634
rect 7657 44582 7669 44634
rect 7669 44582 7699 44634
rect 7723 44582 7733 44634
rect 7733 44582 7779 44634
rect 7483 44580 7539 44582
rect 7563 44580 7619 44582
rect 7643 44580 7699 44582
rect 7723 44580 7779 44582
rect 7483 43546 7539 43548
rect 7563 43546 7619 43548
rect 7643 43546 7699 43548
rect 7723 43546 7779 43548
rect 7483 43494 7529 43546
rect 7529 43494 7539 43546
rect 7563 43494 7593 43546
rect 7593 43494 7605 43546
rect 7605 43494 7619 43546
rect 7643 43494 7657 43546
rect 7657 43494 7669 43546
rect 7669 43494 7699 43546
rect 7723 43494 7733 43546
rect 7733 43494 7779 43546
rect 7483 43492 7539 43494
rect 7563 43492 7619 43494
rect 7643 43492 7699 43494
rect 7723 43492 7779 43494
rect 7483 42458 7539 42460
rect 7563 42458 7619 42460
rect 7643 42458 7699 42460
rect 7723 42458 7779 42460
rect 7483 42406 7529 42458
rect 7529 42406 7539 42458
rect 7563 42406 7593 42458
rect 7593 42406 7605 42458
rect 7605 42406 7619 42458
rect 7643 42406 7657 42458
rect 7657 42406 7669 42458
rect 7669 42406 7699 42458
rect 7723 42406 7733 42458
rect 7733 42406 7779 42458
rect 7483 42404 7539 42406
rect 7563 42404 7619 42406
rect 7643 42404 7699 42406
rect 7723 42404 7779 42406
rect 7483 41370 7539 41372
rect 7563 41370 7619 41372
rect 7643 41370 7699 41372
rect 7723 41370 7779 41372
rect 7483 41318 7529 41370
rect 7529 41318 7539 41370
rect 7563 41318 7593 41370
rect 7593 41318 7605 41370
rect 7605 41318 7619 41370
rect 7643 41318 7657 41370
rect 7657 41318 7669 41370
rect 7669 41318 7699 41370
rect 7723 41318 7733 41370
rect 7733 41318 7779 41370
rect 7483 41316 7539 41318
rect 7563 41316 7619 41318
rect 7643 41316 7699 41318
rect 7723 41316 7779 41318
rect 7483 40282 7539 40284
rect 7563 40282 7619 40284
rect 7643 40282 7699 40284
rect 7723 40282 7779 40284
rect 7483 40230 7529 40282
rect 7529 40230 7539 40282
rect 7563 40230 7593 40282
rect 7593 40230 7605 40282
rect 7605 40230 7619 40282
rect 7643 40230 7657 40282
rect 7657 40230 7669 40282
rect 7669 40230 7699 40282
rect 7723 40230 7733 40282
rect 7733 40230 7779 40282
rect 7483 40228 7539 40230
rect 7563 40228 7619 40230
rect 7643 40228 7699 40230
rect 7723 40228 7779 40230
rect 7483 39194 7539 39196
rect 7563 39194 7619 39196
rect 7643 39194 7699 39196
rect 7723 39194 7779 39196
rect 7483 39142 7529 39194
rect 7529 39142 7539 39194
rect 7563 39142 7593 39194
rect 7593 39142 7605 39194
rect 7605 39142 7619 39194
rect 7643 39142 7657 39194
rect 7657 39142 7669 39194
rect 7669 39142 7699 39194
rect 7723 39142 7733 39194
rect 7733 39142 7779 39194
rect 7483 39140 7539 39142
rect 7563 39140 7619 39142
rect 7643 39140 7699 39142
rect 7723 39140 7779 39142
rect 7483 38106 7539 38108
rect 7563 38106 7619 38108
rect 7643 38106 7699 38108
rect 7723 38106 7779 38108
rect 7483 38054 7529 38106
rect 7529 38054 7539 38106
rect 7563 38054 7593 38106
rect 7593 38054 7605 38106
rect 7605 38054 7619 38106
rect 7643 38054 7657 38106
rect 7657 38054 7669 38106
rect 7669 38054 7699 38106
rect 7723 38054 7733 38106
rect 7733 38054 7779 38106
rect 7483 38052 7539 38054
rect 7563 38052 7619 38054
rect 7643 38052 7699 38054
rect 7723 38052 7779 38054
rect 7483 37018 7539 37020
rect 7563 37018 7619 37020
rect 7643 37018 7699 37020
rect 7723 37018 7779 37020
rect 7483 36966 7529 37018
rect 7529 36966 7539 37018
rect 7563 36966 7593 37018
rect 7593 36966 7605 37018
rect 7605 36966 7619 37018
rect 7643 36966 7657 37018
rect 7657 36966 7669 37018
rect 7669 36966 7699 37018
rect 7723 36966 7733 37018
rect 7733 36966 7779 37018
rect 7483 36964 7539 36966
rect 7563 36964 7619 36966
rect 7643 36964 7699 36966
rect 7723 36964 7779 36966
rect 7483 35930 7539 35932
rect 7563 35930 7619 35932
rect 7643 35930 7699 35932
rect 7723 35930 7779 35932
rect 7483 35878 7529 35930
rect 7529 35878 7539 35930
rect 7563 35878 7593 35930
rect 7593 35878 7605 35930
rect 7605 35878 7619 35930
rect 7643 35878 7657 35930
rect 7657 35878 7669 35930
rect 7669 35878 7699 35930
rect 7723 35878 7733 35930
rect 7733 35878 7779 35930
rect 7483 35876 7539 35878
rect 7563 35876 7619 35878
rect 7643 35876 7699 35878
rect 7723 35876 7779 35878
rect 7483 34842 7539 34844
rect 7563 34842 7619 34844
rect 7643 34842 7699 34844
rect 7723 34842 7779 34844
rect 7483 34790 7529 34842
rect 7529 34790 7539 34842
rect 7563 34790 7593 34842
rect 7593 34790 7605 34842
rect 7605 34790 7619 34842
rect 7643 34790 7657 34842
rect 7657 34790 7669 34842
rect 7669 34790 7699 34842
rect 7723 34790 7733 34842
rect 7733 34790 7779 34842
rect 7483 34788 7539 34790
rect 7563 34788 7619 34790
rect 7643 34788 7699 34790
rect 7723 34788 7779 34790
rect 7483 33754 7539 33756
rect 7563 33754 7619 33756
rect 7643 33754 7699 33756
rect 7723 33754 7779 33756
rect 7483 33702 7529 33754
rect 7529 33702 7539 33754
rect 7563 33702 7593 33754
rect 7593 33702 7605 33754
rect 7605 33702 7619 33754
rect 7643 33702 7657 33754
rect 7657 33702 7669 33754
rect 7669 33702 7699 33754
rect 7723 33702 7733 33754
rect 7733 33702 7779 33754
rect 7483 33700 7539 33702
rect 7563 33700 7619 33702
rect 7643 33700 7699 33702
rect 7723 33700 7779 33702
rect 7483 32666 7539 32668
rect 7563 32666 7619 32668
rect 7643 32666 7699 32668
rect 7723 32666 7779 32668
rect 7483 32614 7529 32666
rect 7529 32614 7539 32666
rect 7563 32614 7593 32666
rect 7593 32614 7605 32666
rect 7605 32614 7619 32666
rect 7643 32614 7657 32666
rect 7657 32614 7669 32666
rect 7669 32614 7699 32666
rect 7723 32614 7733 32666
rect 7733 32614 7779 32666
rect 7483 32612 7539 32614
rect 7563 32612 7619 32614
rect 7643 32612 7699 32614
rect 7723 32612 7779 32614
rect 7483 31578 7539 31580
rect 7563 31578 7619 31580
rect 7643 31578 7699 31580
rect 7723 31578 7779 31580
rect 7483 31526 7529 31578
rect 7529 31526 7539 31578
rect 7563 31526 7593 31578
rect 7593 31526 7605 31578
rect 7605 31526 7619 31578
rect 7643 31526 7657 31578
rect 7657 31526 7669 31578
rect 7669 31526 7699 31578
rect 7723 31526 7733 31578
rect 7733 31526 7779 31578
rect 7483 31524 7539 31526
rect 7563 31524 7619 31526
rect 7643 31524 7699 31526
rect 7723 31524 7779 31526
rect 7483 30490 7539 30492
rect 7563 30490 7619 30492
rect 7643 30490 7699 30492
rect 7723 30490 7779 30492
rect 7483 30438 7529 30490
rect 7529 30438 7539 30490
rect 7563 30438 7593 30490
rect 7593 30438 7605 30490
rect 7605 30438 7619 30490
rect 7643 30438 7657 30490
rect 7657 30438 7669 30490
rect 7669 30438 7699 30490
rect 7723 30438 7733 30490
rect 7733 30438 7779 30490
rect 7483 30436 7539 30438
rect 7563 30436 7619 30438
rect 7643 30436 7699 30438
rect 7723 30436 7779 30438
rect 7483 29402 7539 29404
rect 7563 29402 7619 29404
rect 7643 29402 7699 29404
rect 7723 29402 7779 29404
rect 7483 29350 7529 29402
rect 7529 29350 7539 29402
rect 7563 29350 7593 29402
rect 7593 29350 7605 29402
rect 7605 29350 7619 29402
rect 7643 29350 7657 29402
rect 7657 29350 7669 29402
rect 7669 29350 7699 29402
rect 7723 29350 7733 29402
rect 7733 29350 7779 29402
rect 7483 29348 7539 29350
rect 7563 29348 7619 29350
rect 7643 29348 7699 29350
rect 7723 29348 7779 29350
rect 7483 28314 7539 28316
rect 7563 28314 7619 28316
rect 7643 28314 7699 28316
rect 7723 28314 7779 28316
rect 7483 28262 7529 28314
rect 7529 28262 7539 28314
rect 7563 28262 7593 28314
rect 7593 28262 7605 28314
rect 7605 28262 7619 28314
rect 7643 28262 7657 28314
rect 7657 28262 7669 28314
rect 7669 28262 7699 28314
rect 7723 28262 7733 28314
rect 7733 28262 7779 28314
rect 7483 28260 7539 28262
rect 7563 28260 7619 28262
rect 7643 28260 7699 28262
rect 7723 28260 7779 28262
rect 7483 27226 7539 27228
rect 7563 27226 7619 27228
rect 7643 27226 7699 27228
rect 7723 27226 7779 27228
rect 7483 27174 7529 27226
rect 7529 27174 7539 27226
rect 7563 27174 7593 27226
rect 7593 27174 7605 27226
rect 7605 27174 7619 27226
rect 7643 27174 7657 27226
rect 7657 27174 7669 27226
rect 7669 27174 7699 27226
rect 7723 27174 7733 27226
rect 7733 27174 7779 27226
rect 7483 27172 7539 27174
rect 7563 27172 7619 27174
rect 7643 27172 7699 27174
rect 7723 27172 7779 27174
rect 7483 26138 7539 26140
rect 7563 26138 7619 26140
rect 7643 26138 7699 26140
rect 7723 26138 7779 26140
rect 7483 26086 7529 26138
rect 7529 26086 7539 26138
rect 7563 26086 7593 26138
rect 7593 26086 7605 26138
rect 7605 26086 7619 26138
rect 7643 26086 7657 26138
rect 7657 26086 7669 26138
rect 7669 26086 7699 26138
rect 7723 26086 7733 26138
rect 7733 26086 7779 26138
rect 7483 26084 7539 26086
rect 7563 26084 7619 26086
rect 7643 26084 7699 26086
rect 7723 26084 7779 26086
rect 7483 25050 7539 25052
rect 7563 25050 7619 25052
rect 7643 25050 7699 25052
rect 7723 25050 7779 25052
rect 7483 24998 7529 25050
rect 7529 24998 7539 25050
rect 7563 24998 7593 25050
rect 7593 24998 7605 25050
rect 7605 24998 7619 25050
rect 7643 24998 7657 25050
rect 7657 24998 7669 25050
rect 7669 24998 7699 25050
rect 7723 24998 7733 25050
rect 7733 24998 7779 25050
rect 7483 24996 7539 24998
rect 7563 24996 7619 24998
rect 7643 24996 7699 24998
rect 7723 24996 7779 24998
rect 7483 23962 7539 23964
rect 7563 23962 7619 23964
rect 7643 23962 7699 23964
rect 7723 23962 7779 23964
rect 7483 23910 7529 23962
rect 7529 23910 7539 23962
rect 7563 23910 7593 23962
rect 7593 23910 7605 23962
rect 7605 23910 7619 23962
rect 7643 23910 7657 23962
rect 7657 23910 7669 23962
rect 7669 23910 7699 23962
rect 7723 23910 7733 23962
rect 7733 23910 7779 23962
rect 7483 23908 7539 23910
rect 7563 23908 7619 23910
rect 7643 23908 7699 23910
rect 7723 23908 7779 23910
rect 7483 22874 7539 22876
rect 7563 22874 7619 22876
rect 7643 22874 7699 22876
rect 7723 22874 7779 22876
rect 7483 22822 7529 22874
rect 7529 22822 7539 22874
rect 7563 22822 7593 22874
rect 7593 22822 7605 22874
rect 7605 22822 7619 22874
rect 7643 22822 7657 22874
rect 7657 22822 7669 22874
rect 7669 22822 7699 22874
rect 7723 22822 7733 22874
rect 7733 22822 7779 22874
rect 7483 22820 7539 22822
rect 7563 22820 7619 22822
rect 7643 22820 7699 22822
rect 7723 22820 7779 22822
rect 7483 21786 7539 21788
rect 7563 21786 7619 21788
rect 7643 21786 7699 21788
rect 7723 21786 7779 21788
rect 7483 21734 7529 21786
rect 7529 21734 7539 21786
rect 7563 21734 7593 21786
rect 7593 21734 7605 21786
rect 7605 21734 7619 21786
rect 7643 21734 7657 21786
rect 7657 21734 7669 21786
rect 7669 21734 7699 21786
rect 7723 21734 7733 21786
rect 7733 21734 7779 21786
rect 7483 21732 7539 21734
rect 7563 21732 7619 21734
rect 7643 21732 7699 21734
rect 7723 21732 7779 21734
rect 7483 20698 7539 20700
rect 7563 20698 7619 20700
rect 7643 20698 7699 20700
rect 7723 20698 7779 20700
rect 7483 20646 7529 20698
rect 7529 20646 7539 20698
rect 7563 20646 7593 20698
rect 7593 20646 7605 20698
rect 7605 20646 7619 20698
rect 7643 20646 7657 20698
rect 7657 20646 7669 20698
rect 7669 20646 7699 20698
rect 7723 20646 7733 20698
rect 7733 20646 7779 20698
rect 7483 20644 7539 20646
rect 7563 20644 7619 20646
rect 7643 20644 7699 20646
rect 7723 20644 7779 20646
rect 7483 19610 7539 19612
rect 7563 19610 7619 19612
rect 7643 19610 7699 19612
rect 7723 19610 7779 19612
rect 7483 19558 7529 19610
rect 7529 19558 7539 19610
rect 7563 19558 7593 19610
rect 7593 19558 7605 19610
rect 7605 19558 7619 19610
rect 7643 19558 7657 19610
rect 7657 19558 7669 19610
rect 7669 19558 7699 19610
rect 7723 19558 7733 19610
rect 7733 19558 7779 19610
rect 7483 19556 7539 19558
rect 7563 19556 7619 19558
rect 7643 19556 7699 19558
rect 7723 19556 7779 19558
rect 7483 18522 7539 18524
rect 7563 18522 7619 18524
rect 7643 18522 7699 18524
rect 7723 18522 7779 18524
rect 7483 18470 7529 18522
rect 7529 18470 7539 18522
rect 7563 18470 7593 18522
rect 7593 18470 7605 18522
rect 7605 18470 7619 18522
rect 7643 18470 7657 18522
rect 7657 18470 7669 18522
rect 7669 18470 7699 18522
rect 7723 18470 7733 18522
rect 7733 18470 7779 18522
rect 7483 18468 7539 18470
rect 7563 18468 7619 18470
rect 7643 18468 7699 18470
rect 7723 18468 7779 18470
rect 10046 64368 10102 64424
rect 9115 63674 9171 63676
rect 9195 63674 9251 63676
rect 9275 63674 9331 63676
rect 9355 63674 9411 63676
rect 9115 63622 9161 63674
rect 9161 63622 9171 63674
rect 9195 63622 9225 63674
rect 9225 63622 9237 63674
rect 9237 63622 9251 63674
rect 9275 63622 9289 63674
rect 9289 63622 9301 63674
rect 9301 63622 9331 63674
rect 9355 63622 9365 63674
rect 9365 63622 9411 63674
rect 9115 63620 9171 63622
rect 9195 63620 9251 63622
rect 9275 63620 9331 63622
rect 9355 63620 9411 63622
rect 10046 63552 10102 63608
rect 10046 62872 10102 62928
rect 9115 62586 9171 62588
rect 9195 62586 9251 62588
rect 9275 62586 9331 62588
rect 9355 62586 9411 62588
rect 9115 62534 9161 62586
rect 9161 62534 9171 62586
rect 9195 62534 9225 62586
rect 9225 62534 9237 62586
rect 9237 62534 9251 62586
rect 9275 62534 9289 62586
rect 9289 62534 9301 62586
rect 9301 62534 9331 62586
rect 9355 62534 9365 62586
rect 9365 62534 9411 62586
rect 9115 62532 9171 62534
rect 9195 62532 9251 62534
rect 9275 62532 9331 62534
rect 9355 62532 9411 62534
rect 10046 62092 10048 62112
rect 10048 62092 10100 62112
rect 10100 62092 10102 62112
rect 10046 62056 10102 62092
rect 9115 61498 9171 61500
rect 9195 61498 9251 61500
rect 9275 61498 9331 61500
rect 9355 61498 9411 61500
rect 9115 61446 9161 61498
rect 9161 61446 9171 61498
rect 9195 61446 9225 61498
rect 9225 61446 9237 61498
rect 9237 61446 9251 61498
rect 9275 61446 9289 61498
rect 9289 61446 9301 61498
rect 9301 61446 9331 61498
rect 9355 61446 9365 61498
rect 9365 61446 9411 61498
rect 9115 61444 9171 61446
rect 9195 61444 9251 61446
rect 9275 61444 9331 61446
rect 9355 61444 9411 61446
rect 10046 61376 10102 61432
rect 10046 60580 10102 60616
rect 10046 60560 10048 60580
rect 10048 60560 10100 60580
rect 10100 60560 10102 60580
rect 9115 60410 9171 60412
rect 9195 60410 9251 60412
rect 9275 60410 9331 60412
rect 9355 60410 9411 60412
rect 9115 60358 9161 60410
rect 9161 60358 9171 60410
rect 9195 60358 9225 60410
rect 9225 60358 9237 60410
rect 9237 60358 9251 60410
rect 9275 60358 9289 60410
rect 9289 60358 9301 60410
rect 9301 60358 9331 60410
rect 9355 60358 9365 60410
rect 9365 60358 9411 60410
rect 9115 60356 9171 60358
rect 9195 60356 9251 60358
rect 9275 60356 9331 60358
rect 9355 60356 9411 60358
rect 9115 59322 9171 59324
rect 9195 59322 9251 59324
rect 9275 59322 9331 59324
rect 9355 59322 9411 59324
rect 9115 59270 9161 59322
rect 9161 59270 9171 59322
rect 9195 59270 9225 59322
rect 9225 59270 9237 59322
rect 9237 59270 9251 59322
rect 9275 59270 9289 59322
rect 9289 59270 9301 59322
rect 9301 59270 9331 59322
rect 9355 59270 9365 59322
rect 9365 59270 9411 59322
rect 9115 59268 9171 59270
rect 9195 59268 9251 59270
rect 9275 59268 9331 59270
rect 9355 59268 9411 59270
rect 9115 58234 9171 58236
rect 9195 58234 9251 58236
rect 9275 58234 9331 58236
rect 9355 58234 9411 58236
rect 9115 58182 9161 58234
rect 9161 58182 9171 58234
rect 9195 58182 9225 58234
rect 9225 58182 9237 58234
rect 9237 58182 9251 58234
rect 9275 58182 9289 58234
rect 9289 58182 9301 58234
rect 9301 58182 9331 58234
rect 9355 58182 9365 58234
rect 9365 58182 9411 58234
rect 9115 58180 9171 58182
rect 9195 58180 9251 58182
rect 9275 58180 9331 58182
rect 9355 58180 9411 58182
rect 9115 57146 9171 57148
rect 9195 57146 9251 57148
rect 9275 57146 9331 57148
rect 9355 57146 9411 57148
rect 9115 57094 9161 57146
rect 9161 57094 9171 57146
rect 9195 57094 9225 57146
rect 9225 57094 9237 57146
rect 9237 57094 9251 57146
rect 9275 57094 9289 57146
rect 9289 57094 9301 57146
rect 9301 57094 9331 57146
rect 9355 57094 9365 57146
rect 9365 57094 9411 57146
rect 9115 57092 9171 57094
rect 9195 57092 9251 57094
rect 9275 57092 9331 57094
rect 9355 57092 9411 57094
rect 10046 59916 10048 59936
rect 10048 59916 10100 59936
rect 10100 59916 10102 59936
rect 10046 59880 10102 59916
rect 10046 59064 10102 59120
rect 10046 58404 10102 58440
rect 10046 58384 10048 58404
rect 10048 58384 10100 58404
rect 10100 58384 10102 58404
rect 10046 57568 10102 57624
rect 10046 56888 10102 56944
rect 10046 56108 10048 56128
rect 10048 56108 10100 56128
rect 10100 56108 10102 56128
rect 10046 56072 10102 56108
rect 9115 56058 9171 56060
rect 9195 56058 9251 56060
rect 9275 56058 9331 56060
rect 9355 56058 9411 56060
rect 9115 56006 9161 56058
rect 9161 56006 9171 56058
rect 9195 56006 9225 56058
rect 9225 56006 9237 56058
rect 9237 56006 9251 56058
rect 9275 56006 9289 56058
rect 9289 56006 9301 56058
rect 9301 56006 9331 56058
rect 9355 56006 9365 56058
rect 9365 56006 9411 56058
rect 9115 56004 9171 56006
rect 9195 56004 9251 56006
rect 9275 56004 9331 56006
rect 9355 56004 9411 56006
rect 10046 55256 10102 55312
rect 9115 54970 9171 54972
rect 9195 54970 9251 54972
rect 9275 54970 9331 54972
rect 9355 54970 9411 54972
rect 9115 54918 9161 54970
rect 9161 54918 9171 54970
rect 9195 54918 9225 54970
rect 9225 54918 9237 54970
rect 9237 54918 9251 54970
rect 9275 54918 9289 54970
rect 9289 54918 9301 54970
rect 9301 54918 9331 54970
rect 9355 54918 9365 54970
rect 9365 54918 9411 54970
rect 9115 54916 9171 54918
rect 9195 54916 9251 54918
rect 9275 54916 9331 54918
rect 9355 54916 9411 54918
rect 10138 54612 10140 54632
rect 10140 54612 10192 54632
rect 10192 54612 10194 54632
rect 10138 54576 10194 54612
rect 9115 53882 9171 53884
rect 9195 53882 9251 53884
rect 9275 53882 9331 53884
rect 9355 53882 9411 53884
rect 9115 53830 9161 53882
rect 9161 53830 9171 53882
rect 9195 53830 9225 53882
rect 9225 53830 9237 53882
rect 9237 53830 9251 53882
rect 9275 53830 9289 53882
rect 9289 53830 9301 53882
rect 9301 53830 9331 53882
rect 9355 53830 9365 53882
rect 9365 53830 9411 53882
rect 9115 53828 9171 53830
rect 9195 53828 9251 53830
rect 9275 53828 9331 53830
rect 9355 53828 9411 53830
rect 10138 53760 10194 53816
rect 9115 52794 9171 52796
rect 9195 52794 9251 52796
rect 9275 52794 9331 52796
rect 9355 52794 9411 52796
rect 9115 52742 9161 52794
rect 9161 52742 9171 52794
rect 9195 52742 9225 52794
rect 9225 52742 9237 52794
rect 9237 52742 9251 52794
rect 9275 52742 9289 52794
rect 9289 52742 9301 52794
rect 9301 52742 9331 52794
rect 9355 52742 9365 52794
rect 9365 52742 9411 52794
rect 9115 52740 9171 52742
rect 9195 52740 9251 52742
rect 9275 52740 9331 52742
rect 9355 52740 9411 52742
rect 10138 53080 10194 53136
rect 9115 51706 9171 51708
rect 9195 51706 9251 51708
rect 9275 51706 9331 51708
rect 9355 51706 9411 51708
rect 9115 51654 9161 51706
rect 9161 51654 9171 51706
rect 9195 51654 9225 51706
rect 9225 51654 9237 51706
rect 9237 51654 9251 51706
rect 9275 51654 9289 51706
rect 9289 51654 9301 51706
rect 9301 51654 9331 51706
rect 9355 51654 9365 51706
rect 9365 51654 9411 51706
rect 9115 51652 9171 51654
rect 9195 51652 9251 51654
rect 9275 51652 9331 51654
rect 9355 51652 9411 51654
rect 10138 52264 10194 52320
rect 10138 51584 10194 51640
rect 10138 50768 10194 50824
rect 9115 50618 9171 50620
rect 9195 50618 9251 50620
rect 9275 50618 9331 50620
rect 9355 50618 9411 50620
rect 9115 50566 9161 50618
rect 9161 50566 9171 50618
rect 9195 50566 9225 50618
rect 9225 50566 9237 50618
rect 9237 50566 9251 50618
rect 9275 50566 9289 50618
rect 9289 50566 9301 50618
rect 9301 50566 9331 50618
rect 9355 50566 9365 50618
rect 9365 50566 9411 50618
rect 9115 50564 9171 50566
rect 9195 50564 9251 50566
rect 9275 50564 9331 50566
rect 9355 50564 9411 50566
rect 10138 50088 10194 50144
rect 9115 49530 9171 49532
rect 9195 49530 9251 49532
rect 9275 49530 9331 49532
rect 9355 49530 9411 49532
rect 9115 49478 9161 49530
rect 9161 49478 9171 49530
rect 9195 49478 9225 49530
rect 9225 49478 9237 49530
rect 9237 49478 9251 49530
rect 9275 49478 9289 49530
rect 9289 49478 9301 49530
rect 9301 49478 9331 49530
rect 9355 49478 9365 49530
rect 9365 49478 9411 49530
rect 9115 49476 9171 49478
rect 9195 49476 9251 49478
rect 9275 49476 9331 49478
rect 9355 49476 9411 49478
rect 10138 49272 10194 49328
rect 10138 48592 10194 48648
rect 9115 48442 9171 48444
rect 9195 48442 9251 48444
rect 9275 48442 9331 48444
rect 9355 48442 9411 48444
rect 9115 48390 9161 48442
rect 9161 48390 9171 48442
rect 9195 48390 9225 48442
rect 9225 48390 9237 48442
rect 9237 48390 9251 48442
rect 9275 48390 9289 48442
rect 9289 48390 9301 48442
rect 9301 48390 9331 48442
rect 9355 48390 9365 48442
rect 9365 48390 9411 48442
rect 9115 48388 9171 48390
rect 9195 48388 9251 48390
rect 9275 48388 9331 48390
rect 9355 48388 9411 48390
rect 9115 47354 9171 47356
rect 9195 47354 9251 47356
rect 9275 47354 9331 47356
rect 9355 47354 9411 47356
rect 9115 47302 9161 47354
rect 9161 47302 9171 47354
rect 9195 47302 9225 47354
rect 9225 47302 9237 47354
rect 9237 47302 9251 47354
rect 9275 47302 9289 47354
rect 9289 47302 9301 47354
rect 9301 47302 9331 47354
rect 9355 47302 9365 47354
rect 9365 47302 9411 47354
rect 9115 47300 9171 47302
rect 9195 47300 9251 47302
rect 9275 47300 9331 47302
rect 9355 47300 9411 47302
rect 10138 47776 10194 47832
rect 10138 46996 10140 47016
rect 10140 46996 10192 47016
rect 10192 46996 10194 47016
rect 10138 46960 10194 46996
rect 9115 46266 9171 46268
rect 9195 46266 9251 46268
rect 9275 46266 9331 46268
rect 9355 46266 9411 46268
rect 9115 46214 9161 46266
rect 9161 46214 9171 46266
rect 9195 46214 9225 46266
rect 9225 46214 9237 46266
rect 9237 46214 9251 46266
rect 9275 46214 9289 46266
rect 9289 46214 9301 46266
rect 9301 46214 9331 46266
rect 9355 46214 9365 46266
rect 9365 46214 9411 46266
rect 9115 46212 9171 46214
rect 9195 46212 9251 46214
rect 9275 46212 9331 46214
rect 9355 46212 9411 46214
rect 9115 45178 9171 45180
rect 9195 45178 9251 45180
rect 9275 45178 9331 45180
rect 9355 45178 9411 45180
rect 9115 45126 9161 45178
rect 9161 45126 9171 45178
rect 9195 45126 9225 45178
rect 9225 45126 9237 45178
rect 9237 45126 9251 45178
rect 9275 45126 9289 45178
rect 9289 45126 9301 45178
rect 9301 45126 9331 45178
rect 9355 45126 9365 45178
rect 9365 45126 9411 45178
rect 9115 45124 9171 45126
rect 9195 45124 9251 45126
rect 9275 45124 9331 45126
rect 9355 45124 9411 45126
rect 10138 46280 10194 46336
rect 10138 45464 10194 45520
rect 10138 44820 10140 44840
rect 10140 44820 10192 44840
rect 10192 44820 10194 44840
rect 10138 44784 10194 44820
rect 9115 44090 9171 44092
rect 9195 44090 9251 44092
rect 9275 44090 9331 44092
rect 9355 44090 9411 44092
rect 9115 44038 9161 44090
rect 9161 44038 9171 44090
rect 9195 44038 9225 44090
rect 9225 44038 9237 44090
rect 9237 44038 9251 44090
rect 9275 44038 9289 44090
rect 9289 44038 9301 44090
rect 9301 44038 9331 44090
rect 9355 44038 9365 44090
rect 9365 44038 9411 44090
rect 9115 44036 9171 44038
rect 9195 44036 9251 44038
rect 9275 44036 9331 44038
rect 9355 44036 9411 44038
rect 9115 43002 9171 43004
rect 9195 43002 9251 43004
rect 9275 43002 9331 43004
rect 9355 43002 9411 43004
rect 9115 42950 9161 43002
rect 9161 42950 9171 43002
rect 9195 42950 9225 43002
rect 9225 42950 9237 43002
rect 9237 42950 9251 43002
rect 9275 42950 9289 43002
rect 9289 42950 9301 43002
rect 9301 42950 9331 43002
rect 9355 42950 9365 43002
rect 9365 42950 9411 43002
rect 9115 42948 9171 42950
rect 9195 42948 9251 42950
rect 9275 42948 9331 42950
rect 9355 42948 9411 42950
rect 9115 41914 9171 41916
rect 9195 41914 9251 41916
rect 9275 41914 9331 41916
rect 9355 41914 9411 41916
rect 9115 41862 9161 41914
rect 9161 41862 9171 41914
rect 9195 41862 9225 41914
rect 9225 41862 9237 41914
rect 9237 41862 9251 41914
rect 9275 41862 9289 41914
rect 9289 41862 9301 41914
rect 9301 41862 9331 41914
rect 9355 41862 9365 41914
rect 9365 41862 9411 41914
rect 9115 41860 9171 41862
rect 9195 41860 9251 41862
rect 9275 41860 9331 41862
rect 9355 41860 9411 41862
rect 9115 40826 9171 40828
rect 9195 40826 9251 40828
rect 9275 40826 9331 40828
rect 9355 40826 9411 40828
rect 9115 40774 9161 40826
rect 9161 40774 9171 40826
rect 9195 40774 9225 40826
rect 9225 40774 9237 40826
rect 9237 40774 9251 40826
rect 9275 40774 9289 40826
rect 9289 40774 9301 40826
rect 9301 40774 9331 40826
rect 9355 40774 9365 40826
rect 9365 40774 9411 40826
rect 9115 40772 9171 40774
rect 9195 40772 9251 40774
rect 9275 40772 9331 40774
rect 9355 40772 9411 40774
rect 9115 39738 9171 39740
rect 9195 39738 9251 39740
rect 9275 39738 9331 39740
rect 9355 39738 9411 39740
rect 9115 39686 9161 39738
rect 9161 39686 9171 39738
rect 9195 39686 9225 39738
rect 9225 39686 9237 39738
rect 9237 39686 9251 39738
rect 9275 39686 9289 39738
rect 9289 39686 9301 39738
rect 9301 39686 9331 39738
rect 9355 39686 9365 39738
rect 9365 39686 9411 39738
rect 9115 39684 9171 39686
rect 9195 39684 9251 39686
rect 9275 39684 9331 39686
rect 9355 39684 9411 39686
rect 9115 38650 9171 38652
rect 9195 38650 9251 38652
rect 9275 38650 9331 38652
rect 9355 38650 9411 38652
rect 9115 38598 9161 38650
rect 9161 38598 9171 38650
rect 9195 38598 9225 38650
rect 9225 38598 9237 38650
rect 9237 38598 9251 38650
rect 9275 38598 9289 38650
rect 9289 38598 9301 38650
rect 9301 38598 9331 38650
rect 9355 38598 9365 38650
rect 9365 38598 9411 38650
rect 9115 38596 9171 38598
rect 9195 38596 9251 38598
rect 9275 38596 9331 38598
rect 9355 38596 9411 38598
rect 9115 37562 9171 37564
rect 9195 37562 9251 37564
rect 9275 37562 9331 37564
rect 9355 37562 9411 37564
rect 9115 37510 9161 37562
rect 9161 37510 9171 37562
rect 9195 37510 9225 37562
rect 9225 37510 9237 37562
rect 9237 37510 9251 37562
rect 9275 37510 9289 37562
rect 9289 37510 9301 37562
rect 9301 37510 9331 37562
rect 9355 37510 9365 37562
rect 9365 37510 9411 37562
rect 9115 37508 9171 37510
rect 9195 37508 9251 37510
rect 9275 37508 9331 37510
rect 9355 37508 9411 37510
rect 9115 36474 9171 36476
rect 9195 36474 9251 36476
rect 9275 36474 9331 36476
rect 9355 36474 9411 36476
rect 9115 36422 9161 36474
rect 9161 36422 9171 36474
rect 9195 36422 9225 36474
rect 9225 36422 9237 36474
rect 9237 36422 9251 36474
rect 9275 36422 9289 36474
rect 9289 36422 9301 36474
rect 9301 36422 9331 36474
rect 9355 36422 9365 36474
rect 9365 36422 9411 36474
rect 9115 36420 9171 36422
rect 9195 36420 9251 36422
rect 9275 36420 9331 36422
rect 9355 36420 9411 36422
rect 9115 35386 9171 35388
rect 9195 35386 9251 35388
rect 9275 35386 9331 35388
rect 9355 35386 9411 35388
rect 9115 35334 9161 35386
rect 9161 35334 9171 35386
rect 9195 35334 9225 35386
rect 9225 35334 9237 35386
rect 9237 35334 9251 35386
rect 9275 35334 9289 35386
rect 9289 35334 9301 35386
rect 9301 35334 9331 35386
rect 9355 35334 9365 35386
rect 9365 35334 9411 35386
rect 9115 35332 9171 35334
rect 9195 35332 9251 35334
rect 9275 35332 9331 35334
rect 9355 35332 9411 35334
rect 9115 34298 9171 34300
rect 9195 34298 9251 34300
rect 9275 34298 9331 34300
rect 9355 34298 9411 34300
rect 9115 34246 9161 34298
rect 9161 34246 9171 34298
rect 9195 34246 9225 34298
rect 9225 34246 9237 34298
rect 9237 34246 9251 34298
rect 9275 34246 9289 34298
rect 9289 34246 9301 34298
rect 9301 34246 9331 34298
rect 9355 34246 9365 34298
rect 9365 34246 9411 34298
rect 9115 34244 9171 34246
rect 9195 34244 9251 34246
rect 9275 34244 9331 34246
rect 9355 34244 9411 34246
rect 9115 33210 9171 33212
rect 9195 33210 9251 33212
rect 9275 33210 9331 33212
rect 9355 33210 9411 33212
rect 9115 33158 9161 33210
rect 9161 33158 9171 33210
rect 9195 33158 9225 33210
rect 9225 33158 9237 33210
rect 9237 33158 9251 33210
rect 9275 33158 9289 33210
rect 9289 33158 9301 33210
rect 9301 33158 9331 33210
rect 9355 33158 9365 33210
rect 9365 33158 9411 33210
rect 9115 33156 9171 33158
rect 9195 33156 9251 33158
rect 9275 33156 9331 33158
rect 9355 33156 9411 33158
rect 9115 32122 9171 32124
rect 9195 32122 9251 32124
rect 9275 32122 9331 32124
rect 9355 32122 9411 32124
rect 9115 32070 9161 32122
rect 9161 32070 9171 32122
rect 9195 32070 9225 32122
rect 9225 32070 9237 32122
rect 9237 32070 9251 32122
rect 9275 32070 9289 32122
rect 9289 32070 9301 32122
rect 9301 32070 9331 32122
rect 9355 32070 9365 32122
rect 9365 32070 9411 32122
rect 9115 32068 9171 32070
rect 9195 32068 9251 32070
rect 9275 32068 9331 32070
rect 9355 32068 9411 32070
rect 9115 31034 9171 31036
rect 9195 31034 9251 31036
rect 9275 31034 9331 31036
rect 9355 31034 9411 31036
rect 9115 30982 9161 31034
rect 9161 30982 9171 31034
rect 9195 30982 9225 31034
rect 9225 30982 9237 31034
rect 9237 30982 9251 31034
rect 9275 30982 9289 31034
rect 9289 30982 9301 31034
rect 9301 30982 9331 31034
rect 9355 30982 9365 31034
rect 9365 30982 9411 31034
rect 9115 30980 9171 30982
rect 9195 30980 9251 30982
rect 9275 30980 9331 30982
rect 9355 30980 9411 30982
rect 9115 29946 9171 29948
rect 9195 29946 9251 29948
rect 9275 29946 9331 29948
rect 9355 29946 9411 29948
rect 9115 29894 9161 29946
rect 9161 29894 9171 29946
rect 9195 29894 9225 29946
rect 9225 29894 9237 29946
rect 9237 29894 9251 29946
rect 9275 29894 9289 29946
rect 9289 29894 9301 29946
rect 9301 29894 9331 29946
rect 9355 29894 9365 29946
rect 9365 29894 9411 29946
rect 9115 29892 9171 29894
rect 9195 29892 9251 29894
rect 9275 29892 9331 29894
rect 9355 29892 9411 29894
rect 9115 28858 9171 28860
rect 9195 28858 9251 28860
rect 9275 28858 9331 28860
rect 9355 28858 9411 28860
rect 9115 28806 9161 28858
rect 9161 28806 9171 28858
rect 9195 28806 9225 28858
rect 9225 28806 9237 28858
rect 9237 28806 9251 28858
rect 9275 28806 9289 28858
rect 9289 28806 9301 28858
rect 9301 28806 9331 28858
rect 9355 28806 9365 28858
rect 9365 28806 9411 28858
rect 9115 28804 9171 28806
rect 9195 28804 9251 28806
rect 9275 28804 9331 28806
rect 9355 28804 9411 28806
rect 9115 27770 9171 27772
rect 9195 27770 9251 27772
rect 9275 27770 9331 27772
rect 9355 27770 9411 27772
rect 9115 27718 9161 27770
rect 9161 27718 9171 27770
rect 9195 27718 9225 27770
rect 9225 27718 9237 27770
rect 9237 27718 9251 27770
rect 9275 27718 9289 27770
rect 9289 27718 9301 27770
rect 9301 27718 9331 27770
rect 9355 27718 9365 27770
rect 9365 27718 9411 27770
rect 9115 27716 9171 27718
rect 9195 27716 9251 27718
rect 9275 27716 9331 27718
rect 9355 27716 9411 27718
rect 9115 26682 9171 26684
rect 9195 26682 9251 26684
rect 9275 26682 9331 26684
rect 9355 26682 9411 26684
rect 9115 26630 9161 26682
rect 9161 26630 9171 26682
rect 9195 26630 9225 26682
rect 9225 26630 9237 26682
rect 9237 26630 9251 26682
rect 9275 26630 9289 26682
rect 9289 26630 9301 26682
rect 9301 26630 9331 26682
rect 9355 26630 9365 26682
rect 9365 26630 9411 26682
rect 9115 26628 9171 26630
rect 9195 26628 9251 26630
rect 9275 26628 9331 26630
rect 9355 26628 9411 26630
rect 9115 25594 9171 25596
rect 9195 25594 9251 25596
rect 9275 25594 9331 25596
rect 9355 25594 9411 25596
rect 9115 25542 9161 25594
rect 9161 25542 9171 25594
rect 9195 25542 9225 25594
rect 9225 25542 9237 25594
rect 9237 25542 9251 25594
rect 9275 25542 9289 25594
rect 9289 25542 9301 25594
rect 9301 25542 9331 25594
rect 9355 25542 9365 25594
rect 9365 25542 9411 25594
rect 9115 25540 9171 25542
rect 9195 25540 9251 25542
rect 9275 25540 9331 25542
rect 9355 25540 9411 25542
rect 9115 24506 9171 24508
rect 9195 24506 9251 24508
rect 9275 24506 9331 24508
rect 9355 24506 9411 24508
rect 9115 24454 9161 24506
rect 9161 24454 9171 24506
rect 9195 24454 9225 24506
rect 9225 24454 9237 24506
rect 9237 24454 9251 24506
rect 9275 24454 9289 24506
rect 9289 24454 9301 24506
rect 9301 24454 9331 24506
rect 9355 24454 9365 24506
rect 9365 24454 9411 24506
rect 9115 24452 9171 24454
rect 9195 24452 9251 24454
rect 9275 24452 9331 24454
rect 9355 24452 9411 24454
rect 9115 23418 9171 23420
rect 9195 23418 9251 23420
rect 9275 23418 9331 23420
rect 9355 23418 9411 23420
rect 9115 23366 9161 23418
rect 9161 23366 9171 23418
rect 9195 23366 9225 23418
rect 9225 23366 9237 23418
rect 9237 23366 9251 23418
rect 9275 23366 9289 23418
rect 9289 23366 9301 23418
rect 9301 23366 9331 23418
rect 9355 23366 9365 23418
rect 9365 23366 9411 23418
rect 9115 23364 9171 23366
rect 9195 23364 9251 23366
rect 9275 23364 9331 23366
rect 9355 23364 9411 23366
rect 9126 22888 9182 22944
rect 8850 22072 8906 22128
rect 8942 21392 8998 21448
rect 9115 22330 9171 22332
rect 9195 22330 9251 22332
rect 9275 22330 9331 22332
rect 9355 22330 9411 22332
rect 9115 22278 9161 22330
rect 9161 22278 9171 22330
rect 9195 22278 9225 22330
rect 9225 22278 9237 22330
rect 9237 22278 9251 22330
rect 9275 22278 9289 22330
rect 9289 22278 9301 22330
rect 9301 22278 9331 22330
rect 9355 22278 9365 22330
rect 9365 22278 9411 22330
rect 9115 22276 9171 22278
rect 9195 22276 9251 22278
rect 9275 22276 9331 22278
rect 9355 22276 9411 22278
rect 10138 43968 10194 44024
rect 10138 43288 10194 43344
rect 10138 42472 10194 42528
rect 10138 41792 10194 41848
rect 10138 40976 10194 41032
rect 10138 40296 10194 40352
rect 10138 39480 10194 39536
rect 10138 38664 10194 38720
rect 10138 37984 10194 38040
rect 10138 37204 10140 37224
rect 10140 37204 10192 37224
rect 10192 37204 10194 37224
rect 10138 37168 10194 37204
rect 10138 36488 10194 36544
rect 10138 35672 10194 35728
rect 10138 35028 10140 35048
rect 10140 35028 10192 35048
rect 10192 35028 10194 35048
rect 10138 34992 10194 35028
rect 10138 34176 10194 34232
rect 10138 33496 10194 33552
rect 10138 32680 10194 32736
rect 10138 31864 10194 31920
rect 10138 31184 10194 31240
rect 10138 30368 10194 30424
rect 10138 29688 10194 29744
rect 10138 28872 10194 28928
rect 10138 28192 10194 28248
rect 10138 27376 10194 27432
rect 10230 26696 10286 26752
rect 10046 25880 10102 25936
rect 10138 25236 10140 25256
rect 10140 25236 10192 25256
rect 10192 25236 10194 25256
rect 10138 25200 10194 25236
rect 10138 24384 10194 24440
rect 10138 23568 10194 23624
rect 9115 21242 9171 21244
rect 9195 21242 9251 21244
rect 9275 21242 9331 21244
rect 9355 21242 9411 21244
rect 9115 21190 9161 21242
rect 9161 21190 9171 21242
rect 9195 21190 9225 21242
rect 9225 21190 9237 21242
rect 9237 21190 9251 21242
rect 9275 21190 9289 21242
rect 9289 21190 9301 21242
rect 9301 21190 9331 21242
rect 9355 21190 9365 21242
rect 9365 21190 9411 21242
rect 9115 21188 9171 21190
rect 9195 21188 9251 21190
rect 9275 21188 9331 21190
rect 9355 21188 9411 21190
rect 9034 20576 9090 20632
rect 9115 20154 9171 20156
rect 9195 20154 9251 20156
rect 9275 20154 9331 20156
rect 9355 20154 9411 20156
rect 9115 20102 9161 20154
rect 9161 20102 9171 20154
rect 9195 20102 9225 20154
rect 9225 20102 9237 20154
rect 9237 20102 9251 20154
rect 9275 20102 9289 20154
rect 9289 20102 9301 20154
rect 9301 20102 9331 20154
rect 9355 20102 9365 20154
rect 9365 20102 9411 20154
rect 9115 20100 9171 20102
rect 9195 20100 9251 20102
rect 9275 20100 9331 20102
rect 9355 20100 9411 20102
rect 10138 19896 10194 19952
rect 10230 19080 10286 19136
rect 9115 19066 9171 19068
rect 9195 19066 9251 19068
rect 9275 19066 9331 19068
rect 9355 19066 9411 19068
rect 9115 19014 9161 19066
rect 9161 19014 9171 19066
rect 9195 19014 9225 19066
rect 9225 19014 9237 19066
rect 9237 19014 9251 19066
rect 9275 19014 9289 19066
rect 9289 19014 9301 19066
rect 9301 19014 9331 19066
rect 9355 19014 9365 19066
rect 9365 19014 9411 19066
rect 9115 19012 9171 19014
rect 9195 19012 9251 19014
rect 9275 19012 9331 19014
rect 9355 19012 9411 19014
rect 9115 17978 9171 17980
rect 9195 17978 9251 17980
rect 9275 17978 9331 17980
rect 9355 17978 9411 17980
rect 9115 17926 9161 17978
rect 9161 17926 9171 17978
rect 9195 17926 9225 17978
rect 9225 17926 9237 17978
rect 9237 17926 9251 17978
rect 9275 17926 9289 17978
rect 9289 17926 9301 17978
rect 9301 17926 9331 17978
rect 9355 17926 9365 17978
rect 9365 17926 9411 17978
rect 9115 17924 9171 17926
rect 9195 17924 9251 17926
rect 9275 17924 9331 17926
rect 9355 17924 9411 17926
rect 7483 17434 7539 17436
rect 7563 17434 7619 17436
rect 7643 17434 7699 17436
rect 7723 17434 7779 17436
rect 7483 17382 7529 17434
rect 7529 17382 7539 17434
rect 7563 17382 7593 17434
rect 7593 17382 7605 17434
rect 7605 17382 7619 17434
rect 7643 17382 7657 17434
rect 7657 17382 7669 17434
rect 7669 17382 7699 17434
rect 7723 17382 7733 17434
rect 7733 17382 7779 17434
rect 7483 17380 7539 17382
rect 7563 17380 7619 17382
rect 7643 17380 7699 17382
rect 7723 17380 7779 17382
rect 9115 16890 9171 16892
rect 9195 16890 9251 16892
rect 9275 16890 9331 16892
rect 9355 16890 9411 16892
rect 9115 16838 9161 16890
rect 9161 16838 9171 16890
rect 9195 16838 9225 16890
rect 9225 16838 9237 16890
rect 9237 16838 9251 16890
rect 9275 16838 9289 16890
rect 9289 16838 9301 16890
rect 9301 16838 9331 16890
rect 9355 16838 9365 16890
rect 9365 16838 9411 16890
rect 9115 16836 9171 16838
rect 9195 16836 9251 16838
rect 9275 16836 9331 16838
rect 9355 16836 9411 16838
rect 7483 16346 7539 16348
rect 7563 16346 7619 16348
rect 7643 16346 7699 16348
rect 7723 16346 7779 16348
rect 7483 16294 7529 16346
rect 7529 16294 7539 16346
rect 7563 16294 7593 16346
rect 7593 16294 7605 16346
rect 7605 16294 7619 16346
rect 7643 16294 7657 16346
rect 7657 16294 7669 16346
rect 7669 16294 7699 16346
rect 7723 16294 7733 16346
rect 7733 16294 7779 16346
rect 7483 16292 7539 16294
rect 7563 16292 7619 16294
rect 7643 16292 7699 16294
rect 7723 16292 7779 16294
rect 9115 15802 9171 15804
rect 9195 15802 9251 15804
rect 9275 15802 9331 15804
rect 9355 15802 9411 15804
rect 9115 15750 9161 15802
rect 9161 15750 9171 15802
rect 9195 15750 9225 15802
rect 9225 15750 9237 15802
rect 9237 15750 9251 15802
rect 9275 15750 9289 15802
rect 9289 15750 9301 15802
rect 9301 15750 9331 15802
rect 9355 15750 9365 15802
rect 9365 15750 9411 15802
rect 9115 15748 9171 15750
rect 9195 15748 9251 15750
rect 9275 15748 9331 15750
rect 9355 15748 9411 15750
rect 7483 15258 7539 15260
rect 7563 15258 7619 15260
rect 7643 15258 7699 15260
rect 7723 15258 7779 15260
rect 7483 15206 7529 15258
rect 7529 15206 7539 15258
rect 7563 15206 7593 15258
rect 7593 15206 7605 15258
rect 7605 15206 7619 15258
rect 7643 15206 7657 15258
rect 7657 15206 7669 15258
rect 7669 15206 7699 15258
rect 7723 15206 7733 15258
rect 7733 15206 7779 15258
rect 7483 15204 7539 15206
rect 7563 15204 7619 15206
rect 7643 15204 7699 15206
rect 7723 15204 7779 15206
rect 5851 14714 5907 14716
rect 5931 14714 5987 14716
rect 6011 14714 6067 14716
rect 6091 14714 6147 14716
rect 5851 14662 5897 14714
rect 5897 14662 5907 14714
rect 5931 14662 5961 14714
rect 5961 14662 5973 14714
rect 5973 14662 5987 14714
rect 6011 14662 6025 14714
rect 6025 14662 6037 14714
rect 6037 14662 6067 14714
rect 6091 14662 6101 14714
rect 6101 14662 6147 14714
rect 5851 14660 5907 14662
rect 5931 14660 5987 14662
rect 6011 14660 6067 14662
rect 6091 14660 6147 14662
rect 9115 14714 9171 14716
rect 9195 14714 9251 14716
rect 9275 14714 9331 14716
rect 9355 14714 9411 14716
rect 9115 14662 9161 14714
rect 9161 14662 9171 14714
rect 9195 14662 9225 14714
rect 9225 14662 9237 14714
rect 9237 14662 9251 14714
rect 9275 14662 9289 14714
rect 9289 14662 9301 14714
rect 9301 14662 9331 14714
rect 9355 14662 9365 14714
rect 9365 14662 9411 14714
rect 9115 14660 9171 14662
rect 9195 14660 9251 14662
rect 9275 14660 9331 14662
rect 9355 14660 9411 14662
rect 7483 14170 7539 14172
rect 7563 14170 7619 14172
rect 7643 14170 7699 14172
rect 7723 14170 7779 14172
rect 7483 14118 7529 14170
rect 7529 14118 7539 14170
rect 7563 14118 7593 14170
rect 7593 14118 7605 14170
rect 7605 14118 7619 14170
rect 7643 14118 7657 14170
rect 7657 14118 7669 14170
rect 7669 14118 7699 14170
rect 7723 14118 7733 14170
rect 7733 14118 7779 14170
rect 7483 14116 7539 14118
rect 7563 14116 7619 14118
rect 7643 14116 7699 14118
rect 7723 14116 7779 14118
rect 5851 13626 5907 13628
rect 5931 13626 5987 13628
rect 6011 13626 6067 13628
rect 6091 13626 6147 13628
rect 5851 13574 5897 13626
rect 5897 13574 5907 13626
rect 5931 13574 5961 13626
rect 5961 13574 5973 13626
rect 5973 13574 5987 13626
rect 6011 13574 6025 13626
rect 6025 13574 6037 13626
rect 6037 13574 6067 13626
rect 6091 13574 6101 13626
rect 6101 13574 6147 13626
rect 5851 13572 5907 13574
rect 5931 13572 5987 13574
rect 6011 13572 6067 13574
rect 6091 13572 6147 13574
rect 9115 13626 9171 13628
rect 9195 13626 9251 13628
rect 9275 13626 9331 13628
rect 9355 13626 9411 13628
rect 9115 13574 9161 13626
rect 9161 13574 9171 13626
rect 9195 13574 9225 13626
rect 9225 13574 9237 13626
rect 9237 13574 9251 13626
rect 9275 13574 9289 13626
rect 9289 13574 9301 13626
rect 9301 13574 9331 13626
rect 9355 13574 9365 13626
rect 9365 13574 9411 13626
rect 9115 13572 9171 13574
rect 9195 13572 9251 13574
rect 9275 13572 9331 13574
rect 9355 13572 9411 13574
rect 7483 13082 7539 13084
rect 7563 13082 7619 13084
rect 7643 13082 7699 13084
rect 7723 13082 7779 13084
rect 7483 13030 7529 13082
rect 7529 13030 7539 13082
rect 7563 13030 7593 13082
rect 7593 13030 7605 13082
rect 7605 13030 7619 13082
rect 7643 13030 7657 13082
rect 7657 13030 7669 13082
rect 7669 13030 7699 13082
rect 7723 13030 7733 13082
rect 7733 13030 7779 13082
rect 7483 13028 7539 13030
rect 7563 13028 7619 13030
rect 7643 13028 7699 13030
rect 7723 13028 7779 13030
rect 5851 12538 5907 12540
rect 5931 12538 5987 12540
rect 6011 12538 6067 12540
rect 6091 12538 6147 12540
rect 5851 12486 5897 12538
rect 5897 12486 5907 12538
rect 5931 12486 5961 12538
rect 5961 12486 5973 12538
rect 5973 12486 5987 12538
rect 6011 12486 6025 12538
rect 6025 12486 6037 12538
rect 6037 12486 6067 12538
rect 6091 12486 6101 12538
rect 6101 12486 6147 12538
rect 5851 12484 5907 12486
rect 5931 12484 5987 12486
rect 6011 12484 6067 12486
rect 6091 12484 6147 12486
rect 9115 12538 9171 12540
rect 9195 12538 9251 12540
rect 9275 12538 9331 12540
rect 9355 12538 9411 12540
rect 9115 12486 9161 12538
rect 9161 12486 9171 12538
rect 9195 12486 9225 12538
rect 9225 12486 9237 12538
rect 9237 12486 9251 12538
rect 9275 12486 9289 12538
rect 9289 12486 9301 12538
rect 9301 12486 9331 12538
rect 9355 12486 9365 12538
rect 9365 12486 9411 12538
rect 9115 12484 9171 12486
rect 9195 12484 9251 12486
rect 9275 12484 9331 12486
rect 9355 12484 9411 12486
rect 7483 11994 7539 11996
rect 7563 11994 7619 11996
rect 7643 11994 7699 11996
rect 7723 11994 7779 11996
rect 7483 11942 7529 11994
rect 7529 11942 7539 11994
rect 7563 11942 7593 11994
rect 7593 11942 7605 11994
rect 7605 11942 7619 11994
rect 7643 11942 7657 11994
rect 7657 11942 7669 11994
rect 7669 11942 7699 11994
rect 7723 11942 7733 11994
rect 7733 11942 7779 11994
rect 7483 11940 7539 11942
rect 7563 11940 7619 11942
rect 7643 11940 7699 11942
rect 7723 11940 7779 11942
rect 5851 11450 5907 11452
rect 5931 11450 5987 11452
rect 6011 11450 6067 11452
rect 6091 11450 6147 11452
rect 5851 11398 5897 11450
rect 5897 11398 5907 11450
rect 5931 11398 5961 11450
rect 5961 11398 5973 11450
rect 5973 11398 5987 11450
rect 6011 11398 6025 11450
rect 6025 11398 6037 11450
rect 6037 11398 6067 11450
rect 6091 11398 6101 11450
rect 6101 11398 6147 11450
rect 5851 11396 5907 11398
rect 5931 11396 5987 11398
rect 6011 11396 6067 11398
rect 6091 11396 6147 11398
rect 9115 11450 9171 11452
rect 9195 11450 9251 11452
rect 9275 11450 9331 11452
rect 9355 11450 9411 11452
rect 9115 11398 9161 11450
rect 9161 11398 9171 11450
rect 9195 11398 9225 11450
rect 9225 11398 9237 11450
rect 9237 11398 9251 11450
rect 9275 11398 9289 11450
rect 9289 11398 9301 11450
rect 9301 11398 9331 11450
rect 9355 11398 9365 11450
rect 9365 11398 9411 11450
rect 9115 11396 9171 11398
rect 9195 11396 9251 11398
rect 9275 11396 9331 11398
rect 9355 11396 9411 11398
rect 7483 10906 7539 10908
rect 7563 10906 7619 10908
rect 7643 10906 7699 10908
rect 7723 10906 7779 10908
rect 7483 10854 7529 10906
rect 7529 10854 7539 10906
rect 7563 10854 7593 10906
rect 7593 10854 7605 10906
rect 7605 10854 7619 10906
rect 7643 10854 7657 10906
rect 7657 10854 7669 10906
rect 7669 10854 7699 10906
rect 7723 10854 7733 10906
rect 7733 10854 7779 10906
rect 7483 10852 7539 10854
rect 7563 10852 7619 10854
rect 7643 10852 7699 10854
rect 7723 10852 7779 10854
rect 5851 10362 5907 10364
rect 5931 10362 5987 10364
rect 6011 10362 6067 10364
rect 6091 10362 6147 10364
rect 5851 10310 5897 10362
rect 5897 10310 5907 10362
rect 5931 10310 5961 10362
rect 5961 10310 5973 10362
rect 5973 10310 5987 10362
rect 6011 10310 6025 10362
rect 6025 10310 6037 10362
rect 6037 10310 6067 10362
rect 6091 10310 6101 10362
rect 6101 10310 6147 10362
rect 5851 10308 5907 10310
rect 5931 10308 5987 10310
rect 6011 10308 6067 10310
rect 6091 10308 6147 10310
rect 9115 10362 9171 10364
rect 9195 10362 9251 10364
rect 9275 10362 9331 10364
rect 9355 10362 9411 10364
rect 9115 10310 9161 10362
rect 9161 10310 9171 10362
rect 9195 10310 9225 10362
rect 9225 10310 9237 10362
rect 9237 10310 9251 10362
rect 9275 10310 9289 10362
rect 9289 10310 9301 10362
rect 9301 10310 9331 10362
rect 9355 10310 9365 10362
rect 9365 10310 9411 10362
rect 9115 10308 9171 10310
rect 9195 10308 9251 10310
rect 9275 10308 9331 10310
rect 9355 10308 9411 10310
rect 7483 9818 7539 9820
rect 7563 9818 7619 9820
rect 7643 9818 7699 9820
rect 7723 9818 7779 9820
rect 7483 9766 7529 9818
rect 7529 9766 7539 9818
rect 7563 9766 7593 9818
rect 7593 9766 7605 9818
rect 7605 9766 7619 9818
rect 7643 9766 7657 9818
rect 7657 9766 7669 9818
rect 7669 9766 7699 9818
rect 7723 9766 7733 9818
rect 7733 9766 7779 9818
rect 7483 9764 7539 9766
rect 7563 9764 7619 9766
rect 7643 9764 7699 9766
rect 7723 9764 7779 9766
rect 5851 9274 5907 9276
rect 5931 9274 5987 9276
rect 6011 9274 6067 9276
rect 6091 9274 6147 9276
rect 5851 9222 5897 9274
rect 5897 9222 5907 9274
rect 5931 9222 5961 9274
rect 5961 9222 5973 9274
rect 5973 9222 5987 9274
rect 6011 9222 6025 9274
rect 6025 9222 6037 9274
rect 6037 9222 6067 9274
rect 6091 9222 6101 9274
rect 6101 9222 6147 9274
rect 5851 9220 5907 9222
rect 5931 9220 5987 9222
rect 6011 9220 6067 9222
rect 6091 9220 6147 9222
rect 9115 9274 9171 9276
rect 9195 9274 9251 9276
rect 9275 9274 9331 9276
rect 9355 9274 9411 9276
rect 9115 9222 9161 9274
rect 9161 9222 9171 9274
rect 9195 9222 9225 9274
rect 9225 9222 9237 9274
rect 9237 9222 9251 9274
rect 9275 9222 9289 9274
rect 9289 9222 9301 9274
rect 9301 9222 9331 9274
rect 9355 9222 9365 9274
rect 9365 9222 9411 9274
rect 9115 9220 9171 9222
rect 9195 9220 9251 9222
rect 9275 9220 9331 9222
rect 9355 9220 9411 9222
rect 7483 8730 7539 8732
rect 7563 8730 7619 8732
rect 7643 8730 7699 8732
rect 7723 8730 7779 8732
rect 7483 8678 7529 8730
rect 7529 8678 7539 8730
rect 7563 8678 7593 8730
rect 7593 8678 7605 8730
rect 7605 8678 7619 8730
rect 7643 8678 7657 8730
rect 7657 8678 7669 8730
rect 7669 8678 7699 8730
rect 7723 8678 7733 8730
rect 7733 8678 7779 8730
rect 7483 8676 7539 8678
rect 7563 8676 7619 8678
rect 7643 8676 7699 8678
rect 7723 8676 7779 8678
rect 5851 8186 5907 8188
rect 5931 8186 5987 8188
rect 6011 8186 6067 8188
rect 6091 8186 6147 8188
rect 5851 8134 5897 8186
rect 5897 8134 5907 8186
rect 5931 8134 5961 8186
rect 5961 8134 5973 8186
rect 5973 8134 5987 8186
rect 6011 8134 6025 8186
rect 6025 8134 6037 8186
rect 6037 8134 6067 8186
rect 6091 8134 6101 8186
rect 6101 8134 6147 8186
rect 5851 8132 5907 8134
rect 5931 8132 5987 8134
rect 6011 8132 6067 8134
rect 6091 8132 6147 8134
rect 9115 8186 9171 8188
rect 9195 8186 9251 8188
rect 9275 8186 9331 8188
rect 9355 8186 9411 8188
rect 9115 8134 9161 8186
rect 9161 8134 9171 8186
rect 9195 8134 9225 8186
rect 9225 8134 9237 8186
rect 9237 8134 9251 8186
rect 9275 8134 9289 8186
rect 9289 8134 9301 8186
rect 9301 8134 9331 8186
rect 9355 8134 9365 8186
rect 9365 8134 9411 8186
rect 9115 8132 9171 8134
rect 9195 8132 9251 8134
rect 9275 8132 9331 8134
rect 9355 8132 9411 8134
rect 7483 7642 7539 7644
rect 7563 7642 7619 7644
rect 7643 7642 7699 7644
rect 7723 7642 7779 7644
rect 7483 7590 7529 7642
rect 7529 7590 7539 7642
rect 7563 7590 7593 7642
rect 7593 7590 7605 7642
rect 7605 7590 7619 7642
rect 7643 7590 7657 7642
rect 7657 7590 7669 7642
rect 7669 7590 7699 7642
rect 7723 7590 7733 7642
rect 7733 7590 7779 7642
rect 7483 7588 7539 7590
rect 7563 7588 7619 7590
rect 7643 7588 7699 7590
rect 7723 7588 7779 7590
rect 5851 7098 5907 7100
rect 5931 7098 5987 7100
rect 6011 7098 6067 7100
rect 6091 7098 6147 7100
rect 5851 7046 5897 7098
rect 5897 7046 5907 7098
rect 5931 7046 5961 7098
rect 5961 7046 5973 7098
rect 5973 7046 5987 7098
rect 6011 7046 6025 7098
rect 6025 7046 6037 7098
rect 6037 7046 6067 7098
rect 6091 7046 6101 7098
rect 6101 7046 6147 7098
rect 5851 7044 5907 7046
rect 5931 7044 5987 7046
rect 6011 7044 6067 7046
rect 6091 7044 6147 7046
rect 9115 7098 9171 7100
rect 9195 7098 9251 7100
rect 9275 7098 9331 7100
rect 9355 7098 9411 7100
rect 9115 7046 9161 7098
rect 9161 7046 9171 7098
rect 9195 7046 9225 7098
rect 9225 7046 9237 7098
rect 9237 7046 9251 7098
rect 9275 7046 9289 7098
rect 9289 7046 9301 7098
rect 9301 7046 9331 7098
rect 9355 7046 9365 7098
rect 9365 7046 9411 7098
rect 9115 7044 9171 7046
rect 9195 7044 9251 7046
rect 9275 7044 9331 7046
rect 9355 7044 9411 7046
rect 7483 6554 7539 6556
rect 7563 6554 7619 6556
rect 7643 6554 7699 6556
rect 7723 6554 7779 6556
rect 7483 6502 7529 6554
rect 7529 6502 7539 6554
rect 7563 6502 7593 6554
rect 7593 6502 7605 6554
rect 7605 6502 7619 6554
rect 7643 6502 7657 6554
rect 7657 6502 7669 6554
rect 7669 6502 7699 6554
rect 7723 6502 7733 6554
rect 7733 6502 7779 6554
rect 7483 6500 7539 6502
rect 7563 6500 7619 6502
rect 7643 6500 7699 6502
rect 7723 6500 7779 6502
rect 10138 6296 10194 6352
rect 5851 6010 5907 6012
rect 5931 6010 5987 6012
rect 6011 6010 6067 6012
rect 6091 6010 6147 6012
rect 5851 5958 5897 6010
rect 5897 5958 5907 6010
rect 5931 5958 5961 6010
rect 5961 5958 5973 6010
rect 5973 5958 5987 6010
rect 6011 5958 6025 6010
rect 6025 5958 6037 6010
rect 6037 5958 6067 6010
rect 6091 5958 6101 6010
rect 6101 5958 6147 6010
rect 5851 5956 5907 5958
rect 5931 5956 5987 5958
rect 6011 5956 6067 5958
rect 6091 5956 6147 5958
rect 9115 6010 9171 6012
rect 9195 6010 9251 6012
rect 9275 6010 9331 6012
rect 9355 6010 9411 6012
rect 9115 5958 9161 6010
rect 9161 5958 9171 6010
rect 9195 5958 9225 6010
rect 9225 5958 9237 6010
rect 9237 5958 9251 6010
rect 9275 5958 9289 6010
rect 9289 5958 9301 6010
rect 9301 5958 9331 6010
rect 9355 5958 9365 6010
rect 9365 5958 9411 6010
rect 9115 5956 9171 5958
rect 9195 5956 9251 5958
rect 9275 5956 9331 5958
rect 9355 5956 9411 5958
rect 4219 5466 4275 5468
rect 4299 5466 4355 5468
rect 4379 5466 4435 5468
rect 4459 5466 4515 5468
rect 4219 5414 4265 5466
rect 4265 5414 4275 5466
rect 4299 5414 4329 5466
rect 4329 5414 4341 5466
rect 4341 5414 4355 5466
rect 4379 5414 4393 5466
rect 4393 5414 4405 5466
rect 4405 5414 4435 5466
rect 4459 5414 4469 5466
rect 4469 5414 4515 5466
rect 4219 5412 4275 5414
rect 4299 5412 4355 5414
rect 4379 5412 4435 5414
rect 4459 5412 4515 5414
rect 7483 5466 7539 5468
rect 7563 5466 7619 5468
rect 7643 5466 7699 5468
rect 7723 5466 7779 5468
rect 7483 5414 7529 5466
rect 7529 5414 7539 5466
rect 7563 5414 7593 5466
rect 7593 5414 7605 5466
rect 7605 5414 7619 5466
rect 7643 5414 7657 5466
rect 7657 5414 7669 5466
rect 7669 5414 7699 5466
rect 7723 5414 7733 5466
rect 7733 5414 7779 5466
rect 7483 5412 7539 5414
rect 7563 5412 7619 5414
rect 7643 5412 7699 5414
rect 7723 5412 7779 5414
rect 5851 4922 5907 4924
rect 5931 4922 5987 4924
rect 6011 4922 6067 4924
rect 6091 4922 6147 4924
rect 5851 4870 5897 4922
rect 5897 4870 5907 4922
rect 5931 4870 5961 4922
rect 5961 4870 5973 4922
rect 5973 4870 5987 4922
rect 6011 4870 6025 4922
rect 6025 4870 6037 4922
rect 6037 4870 6067 4922
rect 6091 4870 6101 4922
rect 6101 4870 6147 4922
rect 5851 4868 5907 4870
rect 5931 4868 5987 4870
rect 6011 4868 6067 4870
rect 6091 4868 6147 4870
rect 9115 4922 9171 4924
rect 9195 4922 9251 4924
rect 9275 4922 9331 4924
rect 9355 4922 9411 4924
rect 9115 4870 9161 4922
rect 9161 4870 9171 4922
rect 9195 4870 9225 4922
rect 9225 4870 9237 4922
rect 9237 4870 9251 4922
rect 9275 4870 9289 4922
rect 9289 4870 9301 4922
rect 9301 4870 9331 4922
rect 9355 4870 9365 4922
rect 9365 4870 9411 4922
rect 9115 4868 9171 4870
rect 9195 4868 9251 4870
rect 9275 4868 9331 4870
rect 9355 4868 9411 4870
rect 4219 4378 4275 4380
rect 4299 4378 4355 4380
rect 4379 4378 4435 4380
rect 4459 4378 4515 4380
rect 4219 4326 4265 4378
rect 4265 4326 4275 4378
rect 4299 4326 4329 4378
rect 4329 4326 4341 4378
rect 4341 4326 4355 4378
rect 4379 4326 4393 4378
rect 4393 4326 4405 4378
rect 4405 4326 4435 4378
rect 4459 4326 4469 4378
rect 4469 4326 4515 4378
rect 4219 4324 4275 4326
rect 4299 4324 4355 4326
rect 4379 4324 4435 4326
rect 4459 4324 4515 4326
rect 7483 4378 7539 4380
rect 7563 4378 7619 4380
rect 7643 4378 7699 4380
rect 7723 4378 7779 4380
rect 7483 4326 7529 4378
rect 7529 4326 7539 4378
rect 7563 4326 7593 4378
rect 7593 4326 7605 4378
rect 7605 4326 7619 4378
rect 7643 4326 7657 4378
rect 7657 4326 7669 4378
rect 7669 4326 7699 4378
rect 7723 4326 7733 4378
rect 7733 4326 7779 4378
rect 7483 4324 7539 4326
rect 7563 4324 7619 4326
rect 7643 4324 7699 4326
rect 7723 4324 7779 4326
rect 5851 3834 5907 3836
rect 5931 3834 5987 3836
rect 6011 3834 6067 3836
rect 6091 3834 6147 3836
rect 5851 3782 5897 3834
rect 5897 3782 5907 3834
rect 5931 3782 5961 3834
rect 5961 3782 5973 3834
rect 5973 3782 5987 3834
rect 6011 3782 6025 3834
rect 6025 3782 6037 3834
rect 6037 3782 6067 3834
rect 6091 3782 6101 3834
rect 6101 3782 6147 3834
rect 5851 3780 5907 3782
rect 5931 3780 5987 3782
rect 6011 3780 6067 3782
rect 6091 3780 6147 3782
rect 9115 3834 9171 3836
rect 9195 3834 9251 3836
rect 9275 3834 9331 3836
rect 9355 3834 9411 3836
rect 9115 3782 9161 3834
rect 9161 3782 9171 3834
rect 9195 3782 9225 3834
rect 9225 3782 9237 3834
rect 9237 3782 9251 3834
rect 9275 3782 9289 3834
rect 9289 3782 9301 3834
rect 9301 3782 9331 3834
rect 9355 3782 9365 3834
rect 9365 3782 9411 3834
rect 9115 3780 9171 3782
rect 9195 3780 9251 3782
rect 9275 3780 9331 3782
rect 9355 3780 9411 3782
rect 10138 5480 10194 5536
rect 10138 4800 10194 4856
rect 10138 3984 10194 4040
rect 4219 3290 4275 3292
rect 4299 3290 4355 3292
rect 4379 3290 4435 3292
rect 4459 3290 4515 3292
rect 4219 3238 4265 3290
rect 4265 3238 4275 3290
rect 4299 3238 4329 3290
rect 4329 3238 4341 3290
rect 4341 3238 4355 3290
rect 4379 3238 4393 3290
rect 4393 3238 4405 3290
rect 4405 3238 4435 3290
rect 4459 3238 4469 3290
rect 4469 3238 4515 3290
rect 4219 3236 4275 3238
rect 4299 3236 4355 3238
rect 4379 3236 4435 3238
rect 4459 3236 4515 3238
rect 7483 3290 7539 3292
rect 7563 3290 7619 3292
rect 7643 3290 7699 3292
rect 7723 3290 7779 3292
rect 7483 3238 7529 3290
rect 7529 3238 7539 3290
rect 7563 3238 7593 3290
rect 7593 3238 7605 3290
rect 7605 3238 7619 3290
rect 7643 3238 7657 3290
rect 7657 3238 7669 3290
rect 7669 3238 7699 3290
rect 7723 3238 7733 3290
rect 7733 3238 7779 3290
rect 7483 3236 7539 3238
rect 7563 3236 7619 3238
rect 7643 3236 7699 3238
rect 7723 3236 7779 3238
rect 10138 3304 10194 3360
rect 2588 2746 2644 2748
rect 2668 2746 2724 2748
rect 2748 2746 2804 2748
rect 2828 2746 2884 2748
rect 2588 2694 2634 2746
rect 2634 2694 2644 2746
rect 2668 2694 2698 2746
rect 2698 2694 2710 2746
rect 2710 2694 2724 2746
rect 2748 2694 2762 2746
rect 2762 2694 2774 2746
rect 2774 2694 2804 2746
rect 2828 2694 2838 2746
rect 2838 2694 2884 2746
rect 2588 2692 2644 2694
rect 2668 2692 2724 2694
rect 2748 2692 2804 2694
rect 2828 2692 2884 2694
rect 5851 2746 5907 2748
rect 5931 2746 5987 2748
rect 6011 2746 6067 2748
rect 6091 2746 6147 2748
rect 5851 2694 5897 2746
rect 5897 2694 5907 2746
rect 5931 2694 5961 2746
rect 5961 2694 5973 2746
rect 5973 2694 5987 2746
rect 6011 2694 6025 2746
rect 6025 2694 6037 2746
rect 6037 2694 6067 2746
rect 6091 2694 6101 2746
rect 6101 2694 6147 2746
rect 5851 2692 5907 2694
rect 5931 2692 5987 2694
rect 6011 2692 6067 2694
rect 6091 2692 6147 2694
rect 9115 2746 9171 2748
rect 9195 2746 9251 2748
rect 9275 2746 9331 2748
rect 9355 2746 9411 2748
rect 9115 2694 9161 2746
rect 9161 2694 9171 2746
rect 9195 2694 9225 2746
rect 9225 2694 9237 2746
rect 9237 2694 9251 2746
rect 9275 2694 9289 2746
rect 9289 2694 9301 2746
rect 9301 2694 9331 2746
rect 9355 2694 9365 2746
rect 9365 2694 9411 2746
rect 9115 2692 9171 2694
rect 9195 2692 9251 2694
rect 9275 2692 9331 2694
rect 9355 2692 9411 2694
rect 10138 2488 10194 2544
rect 1490 1944 1546 2000
rect 1398 856 1454 912
rect 4219 2202 4275 2204
rect 4299 2202 4355 2204
rect 4379 2202 4435 2204
rect 4459 2202 4515 2204
rect 4219 2150 4265 2202
rect 4265 2150 4275 2202
rect 4299 2150 4329 2202
rect 4329 2150 4341 2202
rect 4341 2150 4355 2202
rect 4379 2150 4393 2202
rect 4393 2150 4405 2202
rect 4405 2150 4435 2202
rect 4459 2150 4469 2202
rect 4469 2150 4515 2202
rect 4219 2148 4275 2150
rect 4299 2148 4355 2150
rect 4379 2148 4435 2150
rect 4459 2148 4515 2150
rect 7483 2202 7539 2204
rect 7563 2202 7619 2204
rect 7643 2202 7699 2204
rect 7723 2202 7779 2204
rect 7483 2150 7529 2202
rect 7529 2150 7539 2202
rect 7563 2150 7593 2202
rect 7593 2150 7605 2202
rect 7605 2150 7619 2202
rect 7643 2150 7657 2202
rect 7657 2150 7669 2202
rect 7669 2150 7699 2202
rect 7723 2150 7733 2202
rect 7733 2150 7779 2202
rect 7483 2148 7539 2150
rect 7563 2148 7619 2150
rect 7643 2148 7699 2150
rect 7723 2148 7779 2150
rect 10138 1808 10194 1864
rect 3054 1400 3110 1456
rect 2778 312 2834 368
<< metal3 >>
rect 0 79658 800 79688
rect 3785 79658 3851 79661
rect 0 79656 3851 79658
rect 0 79600 3790 79656
rect 3846 79600 3851 79656
rect 0 79598 3851 79600
rect 0 79568 800 79598
rect 3785 79595 3851 79598
rect 9581 79522 9647 79525
rect 11200 79522 12000 79552
rect 9581 79520 12000 79522
rect 9581 79464 9586 79520
rect 9642 79464 12000 79520
rect 9581 79462 12000 79464
rect 9581 79459 9647 79462
rect 11200 79432 12000 79462
rect 0 79114 800 79144
rect 3049 79114 3115 79117
rect 0 79112 3115 79114
rect 0 79056 3054 79112
rect 3110 79056 3115 79112
rect 0 79054 3115 79056
rect 0 79024 800 79054
rect 3049 79051 3115 79054
rect 10961 78706 11027 78709
rect 11200 78706 12000 78736
rect 10961 78704 12000 78706
rect 10961 78648 10966 78704
rect 11022 78648 12000 78704
rect 10961 78646 12000 78648
rect 10961 78643 11027 78646
rect 11200 78616 12000 78646
rect 0 78570 800 78600
rect 1485 78570 1551 78573
rect 0 78568 1551 78570
rect 0 78512 1490 78568
rect 1546 78512 1551 78568
rect 0 78510 1551 78512
rect 0 78480 800 78510
rect 1485 78507 1551 78510
rect 0 78026 800 78056
rect 2957 78026 3023 78029
rect 0 78024 3023 78026
rect 0 77968 2962 78024
rect 3018 77968 3023 78024
rect 0 77966 3023 77968
rect 0 77936 800 77966
rect 2957 77963 3023 77966
rect 9489 78026 9555 78029
rect 11200 78026 12000 78056
rect 9489 78024 12000 78026
rect 9489 77968 9494 78024
rect 9550 77968 12000 78024
rect 9489 77966 12000 77968
rect 9489 77963 9555 77966
rect 11200 77936 12000 77966
rect 2576 77824 2896 77825
rect 2576 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2576 77759 2896 77760
rect 5839 77824 6159 77825
rect 5839 77760 5847 77824
rect 5911 77760 5927 77824
rect 5991 77760 6007 77824
rect 6071 77760 6087 77824
rect 6151 77760 6159 77824
rect 5839 77759 6159 77760
rect 9103 77824 9423 77825
rect 9103 77760 9111 77824
rect 9175 77760 9191 77824
rect 9255 77760 9271 77824
rect 9335 77760 9351 77824
rect 9415 77760 9423 77824
rect 9103 77759 9423 77760
rect 0 77482 800 77512
rect 2037 77482 2103 77485
rect 0 77480 2103 77482
rect 0 77424 2042 77480
rect 2098 77424 2103 77480
rect 0 77422 2103 77424
rect 0 77392 800 77422
rect 2037 77419 2103 77422
rect 4207 77280 4527 77281
rect 4207 77216 4215 77280
rect 4279 77216 4295 77280
rect 4359 77216 4375 77280
rect 4439 77216 4455 77280
rect 4519 77216 4527 77280
rect 4207 77215 4527 77216
rect 7471 77280 7791 77281
rect 7471 77216 7479 77280
rect 7543 77216 7559 77280
rect 7623 77216 7639 77280
rect 7703 77216 7719 77280
rect 7783 77216 7791 77280
rect 7471 77215 7791 77216
rect 10041 77210 10107 77213
rect 11200 77210 12000 77240
rect 10041 77208 12000 77210
rect 10041 77152 10046 77208
rect 10102 77152 12000 77208
rect 10041 77150 12000 77152
rect 10041 77147 10107 77150
rect 11200 77120 12000 77150
rect 0 76938 800 76968
rect 1393 76938 1459 76941
rect 0 76936 1459 76938
rect 0 76880 1398 76936
rect 1454 76880 1459 76936
rect 0 76878 1459 76880
rect 0 76848 800 76878
rect 1393 76875 1459 76878
rect 2576 76736 2896 76737
rect 2576 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2576 76671 2896 76672
rect 5839 76736 6159 76737
rect 5839 76672 5847 76736
rect 5911 76672 5927 76736
rect 5991 76672 6007 76736
rect 6071 76672 6087 76736
rect 6151 76672 6159 76736
rect 5839 76671 6159 76672
rect 9103 76736 9423 76737
rect 9103 76672 9111 76736
rect 9175 76672 9191 76736
rect 9255 76672 9271 76736
rect 9335 76672 9351 76736
rect 9415 76672 9423 76736
rect 9103 76671 9423 76672
rect 10041 76530 10107 76533
rect 11200 76530 12000 76560
rect 10041 76528 12000 76530
rect 10041 76472 10046 76528
rect 10102 76472 12000 76528
rect 10041 76470 12000 76472
rect 10041 76467 10107 76470
rect 11200 76440 12000 76470
rect 0 76394 800 76424
rect 1301 76394 1367 76397
rect 0 76392 1367 76394
rect 0 76336 1306 76392
rect 1362 76336 1367 76392
rect 0 76334 1367 76336
rect 0 76304 800 76334
rect 1301 76331 1367 76334
rect 4207 76192 4527 76193
rect 4207 76128 4215 76192
rect 4279 76128 4295 76192
rect 4359 76128 4375 76192
rect 4439 76128 4455 76192
rect 4519 76128 4527 76192
rect 4207 76127 4527 76128
rect 7471 76192 7791 76193
rect 7471 76128 7479 76192
rect 7543 76128 7559 76192
rect 7623 76128 7639 76192
rect 7703 76128 7719 76192
rect 7783 76128 7791 76192
rect 7471 76127 7791 76128
rect 0 75850 800 75880
rect 1393 75850 1459 75853
rect 0 75848 1459 75850
rect 0 75792 1398 75848
rect 1454 75792 1459 75848
rect 0 75790 1459 75792
rect 0 75760 800 75790
rect 1393 75787 1459 75790
rect 10041 75714 10107 75717
rect 11200 75714 12000 75744
rect 10041 75712 12000 75714
rect 10041 75656 10046 75712
rect 10102 75656 12000 75712
rect 10041 75654 12000 75656
rect 10041 75651 10107 75654
rect 2576 75648 2896 75649
rect 2576 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2576 75583 2896 75584
rect 5839 75648 6159 75649
rect 5839 75584 5847 75648
rect 5911 75584 5927 75648
rect 5991 75584 6007 75648
rect 6071 75584 6087 75648
rect 6151 75584 6159 75648
rect 5839 75583 6159 75584
rect 9103 75648 9423 75649
rect 9103 75584 9111 75648
rect 9175 75584 9191 75648
rect 9255 75584 9271 75648
rect 9335 75584 9351 75648
rect 9415 75584 9423 75648
rect 11200 75624 12000 75654
rect 9103 75583 9423 75584
rect 0 75306 800 75336
rect 2037 75306 2103 75309
rect 0 75304 2103 75306
rect 0 75248 2042 75304
rect 2098 75248 2103 75304
rect 0 75246 2103 75248
rect 0 75216 800 75246
rect 2037 75243 2103 75246
rect 4207 75104 4527 75105
rect 4207 75040 4215 75104
rect 4279 75040 4295 75104
rect 4359 75040 4375 75104
rect 4439 75040 4455 75104
rect 4519 75040 4527 75104
rect 4207 75039 4527 75040
rect 7471 75104 7791 75105
rect 7471 75040 7479 75104
rect 7543 75040 7559 75104
rect 7623 75040 7639 75104
rect 7703 75040 7719 75104
rect 7783 75040 7791 75104
rect 7471 75039 7791 75040
rect 10041 75034 10107 75037
rect 11200 75034 12000 75064
rect 10041 75032 12000 75034
rect 10041 74976 10046 75032
rect 10102 74976 12000 75032
rect 10041 74974 12000 74976
rect 10041 74971 10107 74974
rect 11200 74944 12000 74974
rect 0 74762 800 74792
rect 1301 74762 1367 74765
rect 0 74760 1367 74762
rect 0 74704 1306 74760
rect 1362 74704 1367 74760
rect 0 74702 1367 74704
rect 0 74672 800 74702
rect 1301 74699 1367 74702
rect 2576 74560 2896 74561
rect 2576 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2576 74495 2896 74496
rect 5839 74560 6159 74561
rect 5839 74496 5847 74560
rect 5911 74496 5927 74560
rect 5991 74496 6007 74560
rect 6071 74496 6087 74560
rect 6151 74496 6159 74560
rect 5839 74495 6159 74496
rect 9103 74560 9423 74561
rect 9103 74496 9111 74560
rect 9175 74496 9191 74560
rect 9255 74496 9271 74560
rect 9335 74496 9351 74560
rect 9415 74496 9423 74560
rect 9103 74495 9423 74496
rect 0 74218 800 74248
rect 3785 74218 3851 74221
rect 0 74216 3851 74218
rect 0 74160 3790 74216
rect 3846 74160 3851 74216
rect 0 74158 3851 74160
rect 0 74128 800 74158
rect 3785 74155 3851 74158
rect 10041 74218 10107 74221
rect 11200 74218 12000 74248
rect 10041 74216 12000 74218
rect 10041 74160 10046 74216
rect 10102 74160 12000 74216
rect 10041 74158 12000 74160
rect 10041 74155 10107 74158
rect 11200 74128 12000 74158
rect 4207 74016 4527 74017
rect 4207 73952 4215 74016
rect 4279 73952 4295 74016
rect 4359 73952 4375 74016
rect 4439 73952 4455 74016
rect 4519 73952 4527 74016
rect 4207 73951 4527 73952
rect 7471 74016 7791 74017
rect 7471 73952 7479 74016
rect 7543 73952 7559 74016
rect 7623 73952 7639 74016
rect 7703 73952 7719 74016
rect 7783 73952 7791 74016
rect 7471 73951 7791 73952
rect 0 73674 800 73704
rect 1393 73674 1459 73677
rect 0 73672 1459 73674
rect 0 73616 1398 73672
rect 1454 73616 1459 73672
rect 0 73614 1459 73616
rect 0 73584 800 73614
rect 1393 73611 1459 73614
rect 10041 73538 10107 73541
rect 11200 73538 12000 73568
rect 10041 73536 12000 73538
rect 10041 73480 10046 73536
rect 10102 73480 12000 73536
rect 10041 73478 12000 73480
rect 10041 73475 10107 73478
rect 2576 73472 2896 73473
rect 2576 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2576 73407 2896 73408
rect 5839 73472 6159 73473
rect 5839 73408 5847 73472
rect 5911 73408 5927 73472
rect 5991 73408 6007 73472
rect 6071 73408 6087 73472
rect 6151 73408 6159 73472
rect 5839 73407 6159 73408
rect 9103 73472 9423 73473
rect 9103 73408 9111 73472
rect 9175 73408 9191 73472
rect 9255 73408 9271 73472
rect 9335 73408 9351 73472
rect 9415 73408 9423 73472
rect 11200 73448 12000 73478
rect 9103 73407 9423 73408
rect 0 72994 800 73024
rect 2037 72994 2103 72997
rect 0 72992 2103 72994
rect 0 72936 2042 72992
rect 2098 72936 2103 72992
rect 0 72934 2103 72936
rect 0 72904 800 72934
rect 2037 72931 2103 72934
rect 4207 72928 4527 72929
rect 4207 72864 4215 72928
rect 4279 72864 4295 72928
rect 4359 72864 4375 72928
rect 4439 72864 4455 72928
rect 4519 72864 4527 72928
rect 4207 72863 4527 72864
rect 7471 72928 7791 72929
rect 7471 72864 7479 72928
rect 7543 72864 7559 72928
rect 7623 72864 7639 72928
rect 7703 72864 7719 72928
rect 7783 72864 7791 72928
rect 7471 72863 7791 72864
rect 10041 72722 10107 72725
rect 11200 72722 12000 72752
rect 10041 72720 12000 72722
rect 10041 72664 10046 72720
rect 10102 72664 12000 72720
rect 10041 72662 12000 72664
rect 10041 72659 10107 72662
rect 11200 72632 12000 72662
rect 0 72450 800 72480
rect 1393 72450 1459 72453
rect 0 72448 1459 72450
rect 0 72392 1398 72448
rect 1454 72392 1459 72448
rect 0 72390 1459 72392
rect 0 72360 800 72390
rect 1393 72387 1459 72390
rect 2576 72384 2896 72385
rect 2576 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2576 72319 2896 72320
rect 5839 72384 6159 72385
rect 5839 72320 5847 72384
rect 5911 72320 5927 72384
rect 5991 72320 6007 72384
rect 6071 72320 6087 72384
rect 6151 72320 6159 72384
rect 5839 72319 6159 72320
rect 9103 72384 9423 72385
rect 9103 72320 9111 72384
rect 9175 72320 9191 72384
rect 9255 72320 9271 72384
rect 9335 72320 9351 72384
rect 9415 72320 9423 72384
rect 9103 72319 9423 72320
rect 0 71906 800 71936
rect 1393 71906 1459 71909
rect 0 71904 1459 71906
rect 0 71848 1398 71904
rect 1454 71848 1459 71904
rect 0 71846 1459 71848
rect 0 71816 800 71846
rect 1393 71843 1459 71846
rect 10041 71906 10107 71909
rect 11200 71906 12000 71936
rect 10041 71904 12000 71906
rect 10041 71848 10046 71904
rect 10102 71848 12000 71904
rect 10041 71846 12000 71848
rect 10041 71843 10107 71846
rect 4207 71840 4527 71841
rect 4207 71776 4215 71840
rect 4279 71776 4295 71840
rect 4359 71776 4375 71840
rect 4439 71776 4455 71840
rect 4519 71776 4527 71840
rect 4207 71775 4527 71776
rect 7471 71840 7791 71841
rect 7471 71776 7479 71840
rect 7543 71776 7559 71840
rect 7623 71776 7639 71840
rect 7703 71776 7719 71840
rect 7783 71776 7791 71840
rect 11200 71816 12000 71846
rect 7471 71775 7791 71776
rect 0 71362 800 71392
rect 1393 71362 1459 71365
rect 0 71360 1459 71362
rect 0 71304 1398 71360
rect 1454 71304 1459 71360
rect 0 71302 1459 71304
rect 0 71272 800 71302
rect 1393 71299 1459 71302
rect 2576 71296 2896 71297
rect 2576 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2576 71231 2896 71232
rect 5839 71296 6159 71297
rect 5839 71232 5847 71296
rect 5911 71232 5927 71296
rect 5991 71232 6007 71296
rect 6071 71232 6087 71296
rect 6151 71232 6159 71296
rect 5839 71231 6159 71232
rect 9103 71296 9423 71297
rect 9103 71232 9111 71296
rect 9175 71232 9191 71296
rect 9255 71232 9271 71296
rect 9335 71232 9351 71296
rect 9415 71232 9423 71296
rect 9103 71231 9423 71232
rect 10041 71226 10107 71229
rect 11200 71226 12000 71256
rect 10041 71224 12000 71226
rect 10041 71168 10046 71224
rect 10102 71168 12000 71224
rect 10041 71166 12000 71168
rect 10041 71163 10107 71166
rect 11200 71136 12000 71166
rect 0 70818 800 70848
rect 1393 70818 1459 70821
rect 0 70816 1459 70818
rect 0 70760 1398 70816
rect 1454 70760 1459 70816
rect 0 70758 1459 70760
rect 0 70728 800 70758
rect 1393 70755 1459 70758
rect 4207 70752 4527 70753
rect 4207 70688 4215 70752
rect 4279 70688 4295 70752
rect 4359 70688 4375 70752
rect 4439 70688 4455 70752
rect 4519 70688 4527 70752
rect 4207 70687 4527 70688
rect 7471 70752 7791 70753
rect 7471 70688 7479 70752
rect 7543 70688 7559 70752
rect 7623 70688 7639 70752
rect 7703 70688 7719 70752
rect 7783 70688 7791 70752
rect 7471 70687 7791 70688
rect 10685 70410 10751 70413
rect 11200 70410 12000 70440
rect 10685 70408 12000 70410
rect 10685 70352 10690 70408
rect 10746 70352 12000 70408
rect 10685 70350 12000 70352
rect 10685 70347 10751 70350
rect 11200 70320 12000 70350
rect 0 70274 800 70304
rect 1393 70274 1459 70277
rect 0 70272 1459 70274
rect 0 70216 1398 70272
rect 1454 70216 1459 70272
rect 0 70214 1459 70216
rect 0 70184 800 70214
rect 1393 70211 1459 70214
rect 2576 70208 2896 70209
rect 2576 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2576 70143 2896 70144
rect 5839 70208 6159 70209
rect 5839 70144 5847 70208
rect 5911 70144 5927 70208
rect 5991 70144 6007 70208
rect 6071 70144 6087 70208
rect 6151 70144 6159 70208
rect 5839 70143 6159 70144
rect 9103 70208 9423 70209
rect 9103 70144 9111 70208
rect 9175 70144 9191 70208
rect 9255 70144 9271 70208
rect 9335 70144 9351 70208
rect 9415 70144 9423 70208
rect 9103 70143 9423 70144
rect 0 69730 800 69760
rect 1393 69730 1459 69733
rect 0 69728 1459 69730
rect 0 69672 1398 69728
rect 1454 69672 1459 69728
rect 0 69670 1459 69672
rect 0 69640 800 69670
rect 1393 69667 1459 69670
rect 10041 69730 10107 69733
rect 11200 69730 12000 69760
rect 10041 69728 12000 69730
rect 10041 69672 10046 69728
rect 10102 69672 12000 69728
rect 10041 69670 12000 69672
rect 10041 69667 10107 69670
rect 4207 69664 4527 69665
rect 4207 69600 4215 69664
rect 4279 69600 4295 69664
rect 4359 69600 4375 69664
rect 4439 69600 4455 69664
rect 4519 69600 4527 69664
rect 4207 69599 4527 69600
rect 7471 69664 7791 69665
rect 7471 69600 7479 69664
rect 7543 69600 7559 69664
rect 7623 69600 7639 69664
rect 7703 69600 7719 69664
rect 7783 69600 7791 69664
rect 11200 69640 12000 69670
rect 7471 69599 7791 69600
rect 0 69186 800 69216
rect 1393 69186 1459 69189
rect 0 69184 1459 69186
rect 0 69128 1398 69184
rect 1454 69128 1459 69184
rect 0 69126 1459 69128
rect 0 69096 800 69126
rect 1393 69123 1459 69126
rect 2576 69120 2896 69121
rect 2576 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2576 69055 2896 69056
rect 5839 69120 6159 69121
rect 5839 69056 5847 69120
rect 5911 69056 5927 69120
rect 5991 69056 6007 69120
rect 6071 69056 6087 69120
rect 6151 69056 6159 69120
rect 5839 69055 6159 69056
rect 9103 69120 9423 69121
rect 9103 69056 9111 69120
rect 9175 69056 9191 69120
rect 9255 69056 9271 69120
rect 9335 69056 9351 69120
rect 9415 69056 9423 69120
rect 9103 69055 9423 69056
rect 10041 68914 10107 68917
rect 11200 68914 12000 68944
rect 10041 68912 12000 68914
rect 10041 68856 10046 68912
rect 10102 68856 12000 68912
rect 10041 68854 12000 68856
rect 10041 68851 10107 68854
rect 11200 68824 12000 68854
rect 0 68642 800 68672
rect 1393 68642 1459 68645
rect 0 68640 1459 68642
rect 0 68584 1398 68640
rect 1454 68584 1459 68640
rect 0 68582 1459 68584
rect 0 68552 800 68582
rect 1393 68579 1459 68582
rect 4207 68576 4527 68577
rect 4207 68512 4215 68576
rect 4279 68512 4295 68576
rect 4359 68512 4375 68576
rect 4439 68512 4455 68576
rect 4519 68512 4527 68576
rect 4207 68511 4527 68512
rect 7471 68576 7791 68577
rect 7471 68512 7479 68576
rect 7543 68512 7559 68576
rect 7623 68512 7639 68576
rect 7703 68512 7719 68576
rect 7783 68512 7791 68576
rect 7471 68511 7791 68512
rect 10041 68234 10107 68237
rect 11200 68234 12000 68264
rect 10041 68232 12000 68234
rect 10041 68176 10046 68232
rect 10102 68176 12000 68232
rect 10041 68174 12000 68176
rect 10041 68171 10107 68174
rect 11200 68144 12000 68174
rect 0 68098 800 68128
rect 1393 68098 1459 68101
rect 0 68096 1459 68098
rect 0 68040 1398 68096
rect 1454 68040 1459 68096
rect 0 68038 1459 68040
rect 0 68008 800 68038
rect 1393 68035 1459 68038
rect 2576 68032 2896 68033
rect 2576 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2576 67967 2896 67968
rect 5839 68032 6159 68033
rect 5839 67968 5847 68032
rect 5911 67968 5927 68032
rect 5991 67968 6007 68032
rect 6071 67968 6087 68032
rect 6151 67968 6159 68032
rect 5839 67967 6159 67968
rect 9103 68032 9423 68033
rect 9103 67968 9111 68032
rect 9175 67968 9191 68032
rect 9255 67968 9271 68032
rect 9335 67968 9351 68032
rect 9415 67968 9423 68032
rect 9103 67967 9423 67968
rect 0 67554 800 67584
rect 2221 67554 2287 67557
rect 0 67552 2287 67554
rect 0 67496 2226 67552
rect 2282 67496 2287 67552
rect 0 67494 2287 67496
rect 0 67464 800 67494
rect 2221 67491 2287 67494
rect 4207 67488 4527 67489
rect 4207 67424 4215 67488
rect 4279 67424 4295 67488
rect 4359 67424 4375 67488
rect 4439 67424 4455 67488
rect 4519 67424 4527 67488
rect 4207 67423 4527 67424
rect 7471 67488 7791 67489
rect 7471 67424 7479 67488
rect 7543 67424 7559 67488
rect 7623 67424 7639 67488
rect 7703 67424 7719 67488
rect 7783 67424 7791 67488
rect 7471 67423 7791 67424
rect 10041 67418 10107 67421
rect 11200 67418 12000 67448
rect 10041 67416 12000 67418
rect 10041 67360 10046 67416
rect 10102 67360 12000 67416
rect 10041 67358 12000 67360
rect 10041 67355 10107 67358
rect 11200 67328 12000 67358
rect 0 67010 800 67040
rect 2221 67010 2287 67013
rect 0 67008 2287 67010
rect 0 66952 2226 67008
rect 2282 66952 2287 67008
rect 0 66950 2287 66952
rect 0 66920 800 66950
rect 2221 66947 2287 66950
rect 2576 66944 2896 66945
rect 2576 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2576 66879 2896 66880
rect 5839 66944 6159 66945
rect 5839 66880 5847 66944
rect 5911 66880 5927 66944
rect 5991 66880 6007 66944
rect 6071 66880 6087 66944
rect 6151 66880 6159 66944
rect 5839 66879 6159 66880
rect 9103 66944 9423 66945
rect 9103 66880 9111 66944
rect 9175 66880 9191 66944
rect 9255 66880 9271 66944
rect 9335 66880 9351 66944
rect 9415 66880 9423 66944
rect 9103 66879 9423 66880
rect 10041 66738 10107 66741
rect 11200 66738 12000 66768
rect 10041 66736 12000 66738
rect 10041 66680 10046 66736
rect 10102 66680 12000 66736
rect 10041 66678 12000 66680
rect 10041 66675 10107 66678
rect 11200 66648 12000 66678
rect 3877 66602 3943 66605
rect 3877 66600 3986 66602
rect 3877 66544 3882 66600
rect 3938 66544 3986 66600
rect 3877 66539 3986 66544
rect 0 66330 800 66360
rect 3926 66333 3986 66539
rect 4207 66400 4527 66401
rect 4207 66336 4215 66400
rect 4279 66336 4295 66400
rect 4359 66336 4375 66400
rect 4439 66336 4455 66400
rect 4519 66336 4527 66400
rect 4207 66335 4527 66336
rect 7471 66400 7791 66401
rect 7471 66336 7479 66400
rect 7543 66336 7559 66400
rect 7623 66336 7639 66400
rect 7703 66336 7719 66400
rect 7783 66336 7791 66400
rect 7471 66335 7791 66336
rect 1393 66330 1459 66333
rect 0 66328 1459 66330
rect 0 66272 1398 66328
rect 1454 66272 1459 66328
rect 0 66270 1459 66272
rect 0 66240 800 66270
rect 1393 66267 1459 66270
rect 3877 66328 3986 66333
rect 3877 66272 3882 66328
rect 3938 66272 3986 66328
rect 3877 66270 3986 66272
rect 3877 66267 3943 66270
rect 10041 65922 10107 65925
rect 11200 65922 12000 65952
rect 10041 65920 12000 65922
rect 10041 65864 10046 65920
rect 10102 65864 12000 65920
rect 10041 65862 12000 65864
rect 10041 65859 10107 65862
rect 2576 65856 2896 65857
rect 0 65786 800 65816
rect 2576 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2576 65791 2896 65792
rect 5839 65856 6159 65857
rect 5839 65792 5847 65856
rect 5911 65792 5927 65856
rect 5991 65792 6007 65856
rect 6071 65792 6087 65856
rect 6151 65792 6159 65856
rect 5839 65791 6159 65792
rect 9103 65856 9423 65857
rect 9103 65792 9111 65856
rect 9175 65792 9191 65856
rect 9255 65792 9271 65856
rect 9335 65792 9351 65856
rect 9415 65792 9423 65856
rect 11200 65832 12000 65862
rect 9103 65791 9423 65792
rect 1209 65786 1275 65789
rect 0 65784 1275 65786
rect 0 65728 1214 65784
rect 1270 65728 1275 65784
rect 0 65726 1275 65728
rect 0 65696 800 65726
rect 1209 65723 1275 65726
rect 4207 65312 4527 65313
rect 0 65242 800 65272
rect 4207 65248 4215 65312
rect 4279 65248 4295 65312
rect 4359 65248 4375 65312
rect 4439 65248 4455 65312
rect 4519 65248 4527 65312
rect 4207 65247 4527 65248
rect 7471 65312 7791 65313
rect 7471 65248 7479 65312
rect 7543 65248 7559 65312
rect 7623 65248 7639 65312
rect 7703 65248 7719 65312
rect 7783 65248 7791 65312
rect 7471 65247 7791 65248
rect 1301 65242 1367 65245
rect 0 65240 1367 65242
rect 0 65184 1306 65240
rect 1362 65184 1367 65240
rect 0 65182 1367 65184
rect 0 65152 800 65182
rect 1301 65179 1367 65182
rect 10041 65242 10107 65245
rect 11200 65242 12000 65272
rect 10041 65240 12000 65242
rect 10041 65184 10046 65240
rect 10102 65184 12000 65240
rect 10041 65182 12000 65184
rect 10041 65179 10107 65182
rect 11200 65152 12000 65182
rect 2576 64768 2896 64769
rect 0 64698 800 64728
rect 2576 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2576 64703 2896 64704
rect 5839 64768 6159 64769
rect 5839 64704 5847 64768
rect 5911 64704 5927 64768
rect 5991 64704 6007 64768
rect 6071 64704 6087 64768
rect 6151 64704 6159 64768
rect 5839 64703 6159 64704
rect 9103 64768 9423 64769
rect 9103 64704 9111 64768
rect 9175 64704 9191 64768
rect 9255 64704 9271 64768
rect 9335 64704 9351 64768
rect 9415 64704 9423 64768
rect 9103 64703 9423 64704
rect 1393 64698 1459 64701
rect 0 64696 1459 64698
rect 0 64640 1398 64696
rect 1454 64640 1459 64696
rect 0 64638 1459 64640
rect 0 64608 800 64638
rect 1393 64635 1459 64638
rect 10041 64426 10107 64429
rect 11200 64426 12000 64456
rect 10041 64424 12000 64426
rect 10041 64368 10046 64424
rect 10102 64368 12000 64424
rect 10041 64366 12000 64368
rect 10041 64363 10107 64366
rect 11200 64336 12000 64366
rect 4207 64224 4527 64225
rect 0 64154 800 64184
rect 4207 64160 4215 64224
rect 4279 64160 4295 64224
rect 4359 64160 4375 64224
rect 4439 64160 4455 64224
rect 4519 64160 4527 64224
rect 4207 64159 4527 64160
rect 7471 64224 7791 64225
rect 7471 64160 7479 64224
rect 7543 64160 7559 64224
rect 7623 64160 7639 64224
rect 7703 64160 7719 64224
rect 7783 64160 7791 64224
rect 7471 64159 7791 64160
rect 2773 64154 2839 64157
rect 0 64152 2839 64154
rect 0 64096 2778 64152
rect 2834 64096 2839 64152
rect 0 64094 2839 64096
rect 0 64064 800 64094
rect 2773 64091 2839 64094
rect 1485 64018 1551 64021
rect 2497 64018 2563 64021
rect 1485 64016 2563 64018
rect 1485 63960 1490 64016
rect 1546 63960 2502 64016
rect 2558 63960 2563 64016
rect 1485 63958 2563 63960
rect 1485 63955 1551 63958
rect 2497 63955 2563 63958
rect 2576 63680 2896 63681
rect 0 63610 800 63640
rect 2576 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2576 63615 2896 63616
rect 5839 63680 6159 63681
rect 5839 63616 5847 63680
rect 5911 63616 5927 63680
rect 5991 63616 6007 63680
rect 6071 63616 6087 63680
rect 6151 63616 6159 63680
rect 5839 63615 6159 63616
rect 9103 63680 9423 63681
rect 9103 63616 9111 63680
rect 9175 63616 9191 63680
rect 9255 63616 9271 63680
rect 9335 63616 9351 63680
rect 9415 63616 9423 63680
rect 9103 63615 9423 63616
rect 1301 63610 1367 63613
rect 0 63608 1367 63610
rect 0 63552 1306 63608
rect 1362 63552 1367 63608
rect 0 63550 1367 63552
rect 0 63520 800 63550
rect 1301 63547 1367 63550
rect 10041 63610 10107 63613
rect 11200 63610 12000 63640
rect 10041 63608 12000 63610
rect 10041 63552 10046 63608
rect 10102 63552 12000 63608
rect 10041 63550 12000 63552
rect 10041 63547 10107 63550
rect 11200 63520 12000 63550
rect 4207 63136 4527 63137
rect 0 63066 800 63096
rect 4207 63072 4215 63136
rect 4279 63072 4295 63136
rect 4359 63072 4375 63136
rect 4439 63072 4455 63136
rect 4519 63072 4527 63136
rect 4207 63071 4527 63072
rect 7471 63136 7791 63137
rect 7471 63072 7479 63136
rect 7543 63072 7559 63136
rect 7623 63072 7639 63136
rect 7703 63072 7719 63136
rect 7783 63072 7791 63136
rect 7471 63071 7791 63072
rect 3969 63066 4035 63069
rect 0 63064 4035 63066
rect 0 63008 3974 63064
rect 4030 63008 4035 63064
rect 0 63006 4035 63008
rect 0 62976 800 63006
rect 3969 63003 4035 63006
rect 10041 62930 10107 62933
rect 11200 62930 12000 62960
rect 10041 62928 12000 62930
rect 10041 62872 10046 62928
rect 10102 62872 12000 62928
rect 10041 62870 12000 62872
rect 10041 62867 10107 62870
rect 11200 62840 12000 62870
rect 2773 62794 2839 62797
rect 1396 62792 2839 62794
rect 1396 62736 2778 62792
rect 2834 62736 2839 62792
rect 1396 62734 2839 62736
rect 0 62522 800 62552
rect 1396 62522 1456 62734
rect 2773 62731 2839 62734
rect 2576 62592 2896 62593
rect 2576 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2576 62527 2896 62528
rect 5839 62592 6159 62593
rect 5839 62528 5847 62592
rect 5911 62528 5927 62592
rect 5991 62528 6007 62592
rect 6071 62528 6087 62592
rect 6151 62528 6159 62592
rect 5839 62527 6159 62528
rect 9103 62592 9423 62593
rect 9103 62528 9111 62592
rect 9175 62528 9191 62592
rect 9255 62528 9271 62592
rect 9335 62528 9351 62592
rect 9415 62528 9423 62592
rect 9103 62527 9423 62528
rect 0 62462 1456 62522
rect 0 62432 800 62462
rect 10041 62114 10107 62117
rect 11200 62114 12000 62144
rect 10041 62112 12000 62114
rect 10041 62056 10046 62112
rect 10102 62056 12000 62112
rect 10041 62054 12000 62056
rect 10041 62051 10107 62054
rect 4207 62048 4527 62049
rect 0 61978 800 62008
rect 4207 61984 4215 62048
rect 4279 61984 4295 62048
rect 4359 61984 4375 62048
rect 4439 61984 4455 62048
rect 4519 61984 4527 62048
rect 4207 61983 4527 61984
rect 7471 62048 7791 62049
rect 7471 61984 7479 62048
rect 7543 61984 7559 62048
rect 7623 61984 7639 62048
rect 7703 61984 7719 62048
rect 7783 61984 7791 62048
rect 11200 62024 12000 62054
rect 7471 61983 7791 61984
rect 2313 61978 2379 61981
rect 0 61976 2379 61978
rect 0 61920 2318 61976
rect 2374 61920 2379 61976
rect 0 61918 2379 61920
rect 0 61888 800 61918
rect 2313 61915 2379 61918
rect 2576 61504 2896 61505
rect 0 61434 800 61464
rect 2576 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2576 61439 2896 61440
rect 5839 61504 6159 61505
rect 5839 61440 5847 61504
rect 5911 61440 5927 61504
rect 5991 61440 6007 61504
rect 6071 61440 6087 61504
rect 6151 61440 6159 61504
rect 5839 61439 6159 61440
rect 9103 61504 9423 61505
rect 9103 61440 9111 61504
rect 9175 61440 9191 61504
rect 9255 61440 9271 61504
rect 9335 61440 9351 61504
rect 9415 61440 9423 61504
rect 9103 61439 9423 61440
rect 1485 61434 1551 61437
rect 0 61432 1551 61434
rect 0 61376 1490 61432
rect 1546 61376 1551 61432
rect 0 61374 1551 61376
rect 0 61344 800 61374
rect 1485 61371 1551 61374
rect 10041 61434 10107 61437
rect 11200 61434 12000 61464
rect 10041 61432 12000 61434
rect 10041 61376 10046 61432
rect 10102 61376 12000 61432
rect 10041 61374 12000 61376
rect 10041 61371 10107 61374
rect 11200 61344 12000 61374
rect 4207 60960 4527 60961
rect 0 60890 800 60920
rect 4207 60896 4215 60960
rect 4279 60896 4295 60960
rect 4359 60896 4375 60960
rect 4439 60896 4455 60960
rect 4519 60896 4527 60960
rect 4207 60895 4527 60896
rect 7471 60960 7791 60961
rect 7471 60896 7479 60960
rect 7543 60896 7559 60960
rect 7623 60896 7639 60960
rect 7703 60896 7719 60960
rect 7783 60896 7791 60960
rect 7471 60895 7791 60896
rect 1393 60890 1459 60893
rect 0 60888 1459 60890
rect 0 60832 1398 60888
rect 1454 60832 1459 60888
rect 0 60830 1459 60832
rect 0 60800 800 60830
rect 1393 60827 1459 60830
rect 10041 60618 10107 60621
rect 11200 60618 12000 60648
rect 10041 60616 12000 60618
rect 10041 60560 10046 60616
rect 10102 60560 12000 60616
rect 10041 60558 12000 60560
rect 10041 60555 10107 60558
rect 11200 60528 12000 60558
rect 2576 60416 2896 60417
rect 0 60346 800 60376
rect 2576 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2576 60351 2896 60352
rect 5839 60416 6159 60417
rect 5839 60352 5847 60416
rect 5911 60352 5927 60416
rect 5991 60352 6007 60416
rect 6071 60352 6087 60416
rect 6151 60352 6159 60416
rect 5839 60351 6159 60352
rect 9103 60416 9423 60417
rect 9103 60352 9111 60416
rect 9175 60352 9191 60416
rect 9255 60352 9271 60416
rect 9335 60352 9351 60416
rect 9415 60352 9423 60416
rect 9103 60351 9423 60352
rect 1485 60346 1551 60349
rect 0 60344 1551 60346
rect 0 60288 1490 60344
rect 1546 60288 1551 60344
rect 0 60286 1551 60288
rect 0 60256 800 60286
rect 1485 60283 1551 60286
rect 10041 59938 10107 59941
rect 11200 59938 12000 59968
rect 10041 59936 12000 59938
rect 10041 59880 10046 59936
rect 10102 59880 12000 59936
rect 10041 59878 12000 59880
rect 10041 59875 10107 59878
rect 4207 59872 4527 59873
rect 4207 59808 4215 59872
rect 4279 59808 4295 59872
rect 4359 59808 4375 59872
rect 4439 59808 4455 59872
rect 4519 59808 4527 59872
rect 4207 59807 4527 59808
rect 7471 59872 7791 59873
rect 7471 59808 7479 59872
rect 7543 59808 7559 59872
rect 7623 59808 7639 59872
rect 7703 59808 7719 59872
rect 7783 59808 7791 59872
rect 11200 59848 12000 59878
rect 7471 59807 7791 59808
rect 0 59666 800 59696
rect 1393 59666 1459 59669
rect 0 59664 1459 59666
rect 0 59608 1398 59664
rect 1454 59608 1459 59664
rect 0 59606 1459 59608
rect 0 59576 800 59606
rect 1393 59603 1459 59606
rect 1710 59332 1716 59396
rect 1780 59394 1786 59396
rect 2221 59394 2287 59397
rect 1780 59392 2287 59394
rect 1780 59336 2226 59392
rect 2282 59336 2287 59392
rect 1780 59334 2287 59336
rect 1780 59332 1786 59334
rect 2221 59331 2287 59334
rect 2576 59328 2896 59329
rect 2576 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2576 59263 2896 59264
rect 5839 59328 6159 59329
rect 5839 59264 5847 59328
rect 5911 59264 5927 59328
rect 5991 59264 6007 59328
rect 6071 59264 6087 59328
rect 6151 59264 6159 59328
rect 5839 59263 6159 59264
rect 9103 59328 9423 59329
rect 9103 59264 9111 59328
rect 9175 59264 9191 59328
rect 9255 59264 9271 59328
rect 9335 59264 9351 59328
rect 9415 59264 9423 59328
rect 9103 59263 9423 59264
rect 0 59122 800 59152
rect 1485 59122 1551 59125
rect 0 59120 1551 59122
rect 0 59064 1490 59120
rect 1546 59064 1551 59120
rect 0 59062 1551 59064
rect 0 59032 800 59062
rect 1485 59059 1551 59062
rect 10041 59122 10107 59125
rect 11200 59122 12000 59152
rect 10041 59120 12000 59122
rect 10041 59064 10046 59120
rect 10102 59064 12000 59120
rect 10041 59062 12000 59064
rect 10041 59059 10107 59062
rect 11200 59032 12000 59062
rect 4207 58784 4527 58785
rect 4207 58720 4215 58784
rect 4279 58720 4295 58784
rect 4359 58720 4375 58784
rect 4439 58720 4455 58784
rect 4519 58720 4527 58784
rect 4207 58719 4527 58720
rect 7471 58784 7791 58785
rect 7471 58720 7479 58784
rect 7543 58720 7559 58784
rect 7623 58720 7639 58784
rect 7703 58720 7719 58784
rect 7783 58720 7791 58784
rect 7471 58719 7791 58720
rect 0 58578 800 58608
rect 1393 58578 1459 58581
rect 0 58576 1459 58578
rect 0 58520 1398 58576
rect 1454 58520 1459 58576
rect 0 58518 1459 58520
rect 0 58488 800 58518
rect 1393 58515 1459 58518
rect 10041 58442 10107 58445
rect 11200 58442 12000 58472
rect 10041 58440 12000 58442
rect 10041 58384 10046 58440
rect 10102 58384 12000 58440
rect 10041 58382 12000 58384
rect 10041 58379 10107 58382
rect 11200 58352 12000 58382
rect 2576 58240 2896 58241
rect 2576 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2576 58175 2896 58176
rect 5839 58240 6159 58241
rect 5839 58176 5847 58240
rect 5911 58176 5927 58240
rect 5991 58176 6007 58240
rect 6071 58176 6087 58240
rect 6151 58176 6159 58240
rect 5839 58175 6159 58176
rect 9103 58240 9423 58241
rect 9103 58176 9111 58240
rect 9175 58176 9191 58240
rect 9255 58176 9271 58240
rect 9335 58176 9351 58240
rect 9415 58176 9423 58240
rect 9103 58175 9423 58176
rect 0 58034 800 58064
rect 1485 58034 1551 58037
rect 0 58032 1551 58034
rect 0 57976 1490 58032
rect 1546 57976 1551 58032
rect 0 57974 1551 57976
rect 0 57944 800 57974
rect 1485 57971 1551 57974
rect 1945 57898 2011 57901
rect 1902 57896 2011 57898
rect 1902 57840 1950 57896
rect 2006 57840 2011 57896
rect 1902 57835 2011 57840
rect 1577 57762 1643 57765
rect 1902 57762 1962 57835
rect 1577 57760 1962 57762
rect 1577 57704 1582 57760
rect 1638 57704 1962 57760
rect 1577 57702 1962 57704
rect 1577 57699 1643 57702
rect 4207 57696 4527 57697
rect 4207 57632 4215 57696
rect 4279 57632 4295 57696
rect 4359 57632 4375 57696
rect 4439 57632 4455 57696
rect 4519 57632 4527 57696
rect 4207 57631 4527 57632
rect 7471 57696 7791 57697
rect 7471 57632 7479 57696
rect 7543 57632 7559 57696
rect 7623 57632 7639 57696
rect 7703 57632 7719 57696
rect 7783 57632 7791 57696
rect 7471 57631 7791 57632
rect 10041 57626 10107 57629
rect 11200 57626 12000 57656
rect 10041 57624 12000 57626
rect 10041 57568 10046 57624
rect 10102 57568 12000 57624
rect 10041 57566 12000 57568
rect 10041 57563 10107 57566
rect 11200 57536 12000 57566
rect 0 57490 800 57520
rect 2773 57490 2839 57493
rect 0 57488 2839 57490
rect 0 57432 2778 57488
rect 2834 57432 2839 57488
rect 0 57430 2839 57432
rect 0 57400 800 57430
rect 2773 57427 2839 57430
rect 2576 57152 2896 57153
rect 2576 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2576 57087 2896 57088
rect 5839 57152 6159 57153
rect 5839 57088 5847 57152
rect 5911 57088 5927 57152
rect 5991 57088 6007 57152
rect 6071 57088 6087 57152
rect 6151 57088 6159 57152
rect 5839 57087 6159 57088
rect 9103 57152 9423 57153
rect 9103 57088 9111 57152
rect 9175 57088 9191 57152
rect 9255 57088 9271 57152
rect 9335 57088 9351 57152
rect 9415 57088 9423 57152
rect 9103 57087 9423 57088
rect 0 56946 800 56976
rect 1393 56946 1459 56949
rect 0 56944 1459 56946
rect 0 56888 1398 56944
rect 1454 56888 1459 56944
rect 0 56886 1459 56888
rect 0 56856 800 56886
rect 1393 56883 1459 56886
rect 10041 56946 10107 56949
rect 11200 56946 12000 56976
rect 10041 56944 12000 56946
rect 10041 56888 10046 56944
rect 10102 56888 12000 56944
rect 10041 56886 12000 56888
rect 10041 56883 10107 56886
rect 11200 56856 12000 56886
rect 4207 56608 4527 56609
rect 4207 56544 4215 56608
rect 4279 56544 4295 56608
rect 4359 56544 4375 56608
rect 4439 56544 4455 56608
rect 4519 56544 4527 56608
rect 4207 56543 4527 56544
rect 7471 56608 7791 56609
rect 7471 56544 7479 56608
rect 7543 56544 7559 56608
rect 7623 56544 7639 56608
rect 7703 56544 7719 56608
rect 7783 56544 7791 56608
rect 7471 56543 7791 56544
rect 0 56402 800 56432
rect 3969 56402 4035 56405
rect 0 56400 4035 56402
rect 0 56344 3974 56400
rect 4030 56344 4035 56400
rect 0 56342 4035 56344
rect 0 56312 800 56342
rect 3969 56339 4035 56342
rect 3049 56266 3115 56269
rect 5809 56266 5875 56269
rect 3049 56264 5875 56266
rect 3049 56208 3054 56264
rect 3110 56208 5814 56264
rect 5870 56208 5875 56264
rect 3049 56206 5875 56208
rect 3049 56203 3115 56206
rect 5809 56203 5875 56206
rect 10041 56130 10107 56133
rect 11200 56130 12000 56160
rect 10041 56128 12000 56130
rect 10041 56072 10046 56128
rect 10102 56072 12000 56128
rect 10041 56070 12000 56072
rect 10041 56067 10107 56070
rect 2576 56064 2896 56065
rect 2576 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2576 55999 2896 56000
rect 5839 56064 6159 56065
rect 5839 56000 5847 56064
rect 5911 56000 5927 56064
rect 5991 56000 6007 56064
rect 6071 56000 6087 56064
rect 6151 56000 6159 56064
rect 5839 55999 6159 56000
rect 9103 56064 9423 56065
rect 9103 56000 9111 56064
rect 9175 56000 9191 56064
rect 9255 56000 9271 56064
rect 9335 56000 9351 56064
rect 9415 56000 9423 56064
rect 11200 56040 12000 56070
rect 9103 55999 9423 56000
rect 0 55858 800 55888
rect 2957 55858 3023 55861
rect 0 55856 3023 55858
rect 0 55800 2962 55856
rect 3018 55800 3023 55856
rect 0 55798 3023 55800
rect 0 55768 800 55798
rect 2957 55795 3023 55798
rect 4207 55520 4527 55521
rect 4207 55456 4215 55520
rect 4279 55456 4295 55520
rect 4359 55456 4375 55520
rect 4439 55456 4455 55520
rect 4519 55456 4527 55520
rect 4207 55455 4527 55456
rect 7471 55520 7791 55521
rect 7471 55456 7479 55520
rect 7543 55456 7559 55520
rect 7623 55456 7639 55520
rect 7703 55456 7719 55520
rect 7783 55456 7791 55520
rect 7471 55455 7791 55456
rect 0 55314 800 55344
rect 3969 55314 4035 55317
rect 0 55312 4035 55314
rect 0 55256 3974 55312
rect 4030 55256 4035 55312
rect 0 55254 4035 55256
rect 0 55224 800 55254
rect 3969 55251 4035 55254
rect 10041 55314 10107 55317
rect 11200 55314 12000 55344
rect 10041 55312 12000 55314
rect 10041 55256 10046 55312
rect 10102 55256 12000 55312
rect 10041 55254 12000 55256
rect 10041 55251 10107 55254
rect 11200 55224 12000 55254
rect 2576 54976 2896 54977
rect 2576 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2576 54911 2896 54912
rect 5839 54976 6159 54977
rect 5839 54912 5847 54976
rect 5911 54912 5927 54976
rect 5991 54912 6007 54976
rect 6071 54912 6087 54976
rect 6151 54912 6159 54976
rect 5839 54911 6159 54912
rect 9103 54976 9423 54977
rect 9103 54912 9111 54976
rect 9175 54912 9191 54976
rect 9255 54912 9271 54976
rect 9335 54912 9351 54976
rect 9415 54912 9423 54976
rect 9103 54911 9423 54912
rect 0 54770 800 54800
rect 2957 54770 3023 54773
rect 0 54768 3023 54770
rect 0 54712 2962 54768
rect 3018 54712 3023 54768
rect 0 54710 3023 54712
rect 0 54680 800 54710
rect 2957 54707 3023 54710
rect 10133 54634 10199 54637
rect 11200 54634 12000 54664
rect 10133 54632 12000 54634
rect 10133 54576 10138 54632
rect 10194 54576 12000 54632
rect 10133 54574 12000 54576
rect 10133 54571 10199 54574
rect 11200 54544 12000 54574
rect 4207 54432 4527 54433
rect 4207 54368 4215 54432
rect 4279 54368 4295 54432
rect 4359 54368 4375 54432
rect 4439 54368 4455 54432
rect 4519 54368 4527 54432
rect 4207 54367 4527 54368
rect 7471 54432 7791 54433
rect 7471 54368 7479 54432
rect 7543 54368 7559 54432
rect 7623 54368 7639 54432
rect 7703 54368 7719 54432
rect 7783 54368 7791 54432
rect 7471 54367 7791 54368
rect 0 54226 800 54256
rect 1485 54226 1551 54229
rect 0 54224 1551 54226
rect 0 54168 1490 54224
rect 1546 54168 1551 54224
rect 0 54166 1551 54168
rect 0 54136 800 54166
rect 1485 54163 1551 54166
rect 2576 53888 2896 53889
rect 2576 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2576 53823 2896 53824
rect 5839 53888 6159 53889
rect 5839 53824 5847 53888
rect 5911 53824 5927 53888
rect 5991 53824 6007 53888
rect 6071 53824 6087 53888
rect 6151 53824 6159 53888
rect 5839 53823 6159 53824
rect 9103 53888 9423 53889
rect 9103 53824 9111 53888
rect 9175 53824 9191 53888
rect 9255 53824 9271 53888
rect 9335 53824 9351 53888
rect 9415 53824 9423 53888
rect 9103 53823 9423 53824
rect 10133 53818 10199 53821
rect 11200 53818 12000 53848
rect 10133 53816 12000 53818
rect 10133 53760 10138 53816
rect 10194 53760 12000 53816
rect 10133 53758 12000 53760
rect 10133 53755 10199 53758
rect 11200 53728 12000 53758
rect 0 53682 800 53712
rect 1485 53682 1551 53685
rect 0 53680 1551 53682
rect 0 53624 1490 53680
rect 1546 53624 1551 53680
rect 0 53622 1551 53624
rect 0 53592 800 53622
rect 1485 53619 1551 53622
rect 4207 53344 4527 53345
rect 4207 53280 4215 53344
rect 4279 53280 4295 53344
rect 4359 53280 4375 53344
rect 4439 53280 4455 53344
rect 4519 53280 4527 53344
rect 4207 53279 4527 53280
rect 7471 53344 7791 53345
rect 7471 53280 7479 53344
rect 7543 53280 7559 53344
rect 7623 53280 7639 53344
rect 7703 53280 7719 53344
rect 7783 53280 7791 53344
rect 7471 53279 7791 53280
rect 3233 53138 3299 53141
rect 10133 53138 10199 53141
rect 11200 53138 12000 53168
rect 3233 53136 3572 53138
rect 3233 53080 3238 53136
rect 3294 53080 3572 53136
rect 3233 53078 3572 53080
rect 3233 53075 3299 53078
rect 0 53002 800 53032
rect 1485 53002 1551 53005
rect 0 53000 1551 53002
rect 0 52944 1490 53000
rect 1546 52944 1551 53000
rect 0 52942 1551 52944
rect 0 52912 800 52942
rect 1485 52939 1551 52942
rect 2773 53002 2839 53005
rect 2773 53000 3020 53002
rect 2773 52944 2778 53000
rect 2834 52944 3020 53000
rect 2773 52942 3020 52944
rect 2773 52939 2839 52942
rect 2960 52866 3020 52942
rect 3141 52866 3207 52869
rect 2960 52864 3207 52866
rect 2960 52808 3146 52864
rect 3202 52808 3207 52864
rect 2960 52806 3207 52808
rect 3141 52803 3207 52806
rect 2576 52800 2896 52801
rect 2576 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2576 52735 2896 52736
rect 0 52458 800 52488
rect 1485 52458 1551 52461
rect 0 52456 1551 52458
rect 0 52400 1490 52456
rect 1546 52400 1551 52456
rect 0 52398 1551 52400
rect 0 52368 800 52398
rect 1485 52395 1551 52398
rect 3512 52325 3572 53078
rect 10133 53136 12000 53138
rect 10133 53080 10138 53136
rect 10194 53080 12000 53136
rect 10133 53078 12000 53080
rect 10133 53075 10199 53078
rect 11200 53048 12000 53078
rect 5839 52800 6159 52801
rect 5839 52736 5847 52800
rect 5911 52736 5927 52800
rect 5991 52736 6007 52800
rect 6071 52736 6087 52800
rect 6151 52736 6159 52800
rect 5839 52735 6159 52736
rect 9103 52800 9423 52801
rect 9103 52736 9111 52800
rect 9175 52736 9191 52800
rect 9255 52736 9271 52800
rect 9335 52736 9351 52800
rect 9415 52736 9423 52800
rect 9103 52735 9423 52736
rect 3509 52320 3575 52325
rect 3509 52264 3514 52320
rect 3570 52264 3575 52320
rect 3509 52259 3575 52264
rect 10133 52322 10199 52325
rect 11200 52322 12000 52352
rect 10133 52320 12000 52322
rect 10133 52264 10138 52320
rect 10194 52264 12000 52320
rect 10133 52262 12000 52264
rect 10133 52259 10199 52262
rect 4207 52256 4527 52257
rect 4207 52192 4215 52256
rect 4279 52192 4295 52256
rect 4359 52192 4375 52256
rect 4439 52192 4455 52256
rect 4519 52192 4527 52256
rect 4207 52191 4527 52192
rect 7471 52256 7791 52257
rect 7471 52192 7479 52256
rect 7543 52192 7559 52256
rect 7623 52192 7639 52256
rect 7703 52192 7719 52256
rect 7783 52192 7791 52256
rect 11200 52232 12000 52262
rect 7471 52191 7791 52192
rect 2497 52186 2563 52189
rect 3233 52186 3299 52189
rect 2497 52184 3299 52186
rect 2497 52128 2502 52184
rect 2558 52128 3238 52184
rect 3294 52128 3299 52184
rect 2497 52126 3299 52128
rect 2497 52123 2563 52126
rect 3233 52123 3299 52126
rect 0 51914 800 51944
rect 2773 51914 2839 51917
rect 0 51912 2839 51914
rect 0 51856 2778 51912
rect 2834 51856 2839 51912
rect 0 51854 2839 51856
rect 0 51824 800 51854
rect 2773 51851 2839 51854
rect 2576 51712 2896 51713
rect 2576 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2576 51647 2896 51648
rect 5839 51712 6159 51713
rect 5839 51648 5847 51712
rect 5911 51648 5927 51712
rect 5991 51648 6007 51712
rect 6071 51648 6087 51712
rect 6151 51648 6159 51712
rect 5839 51647 6159 51648
rect 9103 51712 9423 51713
rect 9103 51648 9111 51712
rect 9175 51648 9191 51712
rect 9255 51648 9271 51712
rect 9335 51648 9351 51712
rect 9415 51648 9423 51712
rect 9103 51647 9423 51648
rect 2313 51642 2379 51645
rect 2270 51640 2379 51642
rect 2270 51584 2318 51640
rect 2374 51584 2379 51640
rect 2270 51579 2379 51584
rect 10133 51642 10199 51645
rect 11200 51642 12000 51672
rect 10133 51640 12000 51642
rect 10133 51584 10138 51640
rect 10194 51584 12000 51640
rect 10133 51582 12000 51584
rect 10133 51579 10199 51582
rect 0 51370 800 51400
rect 1485 51370 1551 51373
rect 0 51368 1551 51370
rect 0 51312 1490 51368
rect 1546 51312 1551 51368
rect 0 51310 1551 51312
rect 0 51280 800 51310
rect 1485 51307 1551 51310
rect 2270 51101 2330 51579
rect 11200 51552 12000 51582
rect 2405 51506 2471 51509
rect 7833 51506 7899 51509
rect 2405 51504 7899 51506
rect 2405 51448 2410 51504
rect 2466 51448 7838 51504
rect 7894 51448 7899 51504
rect 2405 51446 7899 51448
rect 2405 51443 2471 51446
rect 7833 51443 7899 51446
rect 2589 51370 2655 51373
rect 5809 51370 5875 51373
rect 2589 51368 5875 51370
rect 2589 51312 2594 51368
rect 2650 51312 5814 51368
rect 5870 51312 5875 51368
rect 2589 51310 5875 51312
rect 2589 51307 2655 51310
rect 5809 51307 5875 51310
rect 4207 51168 4527 51169
rect 4207 51104 4215 51168
rect 4279 51104 4295 51168
rect 4359 51104 4375 51168
rect 4439 51104 4455 51168
rect 4519 51104 4527 51168
rect 4207 51103 4527 51104
rect 7471 51168 7791 51169
rect 7471 51104 7479 51168
rect 7543 51104 7559 51168
rect 7623 51104 7639 51168
rect 7703 51104 7719 51168
rect 7783 51104 7791 51168
rect 7471 51103 7791 51104
rect 2221 51096 2330 51101
rect 2221 51040 2226 51096
rect 2282 51040 2330 51096
rect 2221 51038 2330 51040
rect 3969 51088 4035 51093
rect 2221 51035 2287 51038
rect 3969 51032 3974 51088
rect 4030 51032 4035 51088
rect 3969 51027 4035 51032
rect 1669 50964 1735 50965
rect 1669 50960 1716 50964
rect 1780 50962 1786 50964
rect 3972 50962 4032 51027
rect 1669 50904 1674 50960
rect 1669 50900 1716 50904
rect 1780 50902 1826 50962
rect 3926 50902 4032 50962
rect 1780 50900 1786 50902
rect 1669 50899 1735 50900
rect 0 50826 800 50856
rect 2773 50826 2839 50829
rect 0 50824 2839 50826
rect 0 50768 2778 50824
rect 2834 50768 2839 50824
rect 0 50766 2839 50768
rect 0 50736 800 50766
rect 2773 50763 2839 50766
rect 3509 50826 3575 50829
rect 3926 50826 3986 50902
rect 3509 50824 3986 50826
rect 3509 50768 3514 50824
rect 3570 50768 3986 50824
rect 3509 50766 3986 50768
rect 10133 50826 10199 50829
rect 11200 50826 12000 50856
rect 10133 50824 12000 50826
rect 10133 50768 10138 50824
rect 10194 50768 12000 50824
rect 10133 50766 12000 50768
rect 3509 50763 3575 50766
rect 10133 50763 10199 50766
rect 11200 50736 12000 50766
rect 2576 50624 2896 50625
rect 2576 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2576 50559 2896 50560
rect 5839 50624 6159 50625
rect 5839 50560 5847 50624
rect 5911 50560 5927 50624
rect 5991 50560 6007 50624
rect 6071 50560 6087 50624
rect 6151 50560 6159 50624
rect 5839 50559 6159 50560
rect 9103 50624 9423 50625
rect 9103 50560 9111 50624
rect 9175 50560 9191 50624
rect 9255 50560 9271 50624
rect 9335 50560 9351 50624
rect 9415 50560 9423 50624
rect 9103 50559 9423 50560
rect 0 50282 800 50312
rect 2497 50282 2563 50285
rect 0 50280 2563 50282
rect 0 50224 2502 50280
rect 2558 50224 2563 50280
rect 0 50222 2563 50224
rect 0 50192 800 50222
rect 2497 50219 2563 50222
rect 10133 50146 10199 50149
rect 11200 50146 12000 50176
rect 10133 50144 12000 50146
rect 10133 50088 10138 50144
rect 10194 50088 12000 50144
rect 10133 50086 12000 50088
rect 10133 50083 10199 50086
rect 4207 50080 4527 50081
rect 4207 50016 4215 50080
rect 4279 50016 4295 50080
rect 4359 50016 4375 50080
rect 4439 50016 4455 50080
rect 4519 50016 4527 50080
rect 4207 50015 4527 50016
rect 7471 50080 7791 50081
rect 7471 50016 7479 50080
rect 7543 50016 7559 50080
rect 7623 50016 7639 50080
rect 7703 50016 7719 50080
rect 7783 50016 7791 50080
rect 11200 50056 12000 50086
rect 7471 50015 7791 50016
rect 0 49738 800 49768
rect 1485 49738 1551 49741
rect 0 49736 1551 49738
rect 0 49680 1490 49736
rect 1546 49680 1551 49736
rect 0 49678 1551 49680
rect 0 49648 800 49678
rect 1485 49675 1551 49678
rect 2576 49536 2896 49537
rect 2576 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2576 49471 2896 49472
rect 5839 49536 6159 49537
rect 5839 49472 5847 49536
rect 5911 49472 5927 49536
rect 5991 49472 6007 49536
rect 6071 49472 6087 49536
rect 6151 49472 6159 49536
rect 5839 49471 6159 49472
rect 9103 49536 9423 49537
rect 9103 49472 9111 49536
rect 9175 49472 9191 49536
rect 9255 49472 9271 49536
rect 9335 49472 9351 49536
rect 9415 49472 9423 49536
rect 9103 49471 9423 49472
rect 10133 49330 10199 49333
rect 11200 49330 12000 49360
rect 10133 49328 12000 49330
rect 10133 49272 10138 49328
rect 10194 49272 12000 49328
rect 10133 49270 12000 49272
rect 10133 49267 10199 49270
rect 11200 49240 12000 49270
rect 0 49194 800 49224
rect 1485 49194 1551 49197
rect 0 49192 1551 49194
rect 0 49136 1490 49192
rect 1546 49136 1551 49192
rect 0 49134 1551 49136
rect 0 49104 800 49134
rect 1485 49131 1551 49134
rect 4207 48992 4527 48993
rect 4207 48928 4215 48992
rect 4279 48928 4295 48992
rect 4359 48928 4375 48992
rect 4439 48928 4455 48992
rect 4519 48928 4527 48992
rect 4207 48927 4527 48928
rect 7471 48992 7791 48993
rect 7471 48928 7479 48992
rect 7543 48928 7559 48992
rect 7623 48928 7639 48992
rect 7703 48928 7719 48992
rect 7783 48928 7791 48992
rect 7471 48927 7791 48928
rect 0 48650 800 48680
rect 1485 48650 1551 48653
rect 0 48648 1551 48650
rect 0 48592 1490 48648
rect 1546 48592 1551 48648
rect 0 48590 1551 48592
rect 0 48560 800 48590
rect 1485 48587 1551 48590
rect 3693 48650 3759 48653
rect 10133 48650 10199 48653
rect 11200 48650 12000 48680
rect 3693 48648 3802 48650
rect 3693 48592 3698 48648
rect 3754 48592 3802 48648
rect 3693 48587 3802 48592
rect 10133 48648 12000 48650
rect 10133 48592 10138 48648
rect 10194 48592 12000 48648
rect 10133 48590 12000 48592
rect 10133 48587 10199 48590
rect 2576 48448 2896 48449
rect 2576 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2576 48383 2896 48384
rect 3742 48381 3802 48587
rect 11200 48560 12000 48590
rect 5839 48448 6159 48449
rect 5839 48384 5847 48448
rect 5911 48384 5927 48448
rect 5991 48384 6007 48448
rect 6071 48384 6087 48448
rect 6151 48384 6159 48448
rect 5839 48383 6159 48384
rect 9103 48448 9423 48449
rect 9103 48384 9111 48448
rect 9175 48384 9191 48448
rect 9255 48384 9271 48448
rect 9335 48384 9351 48448
rect 9415 48384 9423 48448
rect 9103 48383 9423 48384
rect 3693 48376 3802 48381
rect 3693 48320 3698 48376
rect 3754 48320 3802 48376
rect 3693 48318 3802 48320
rect 3693 48315 3759 48318
rect 0 48106 800 48136
rect 1485 48106 1551 48109
rect 0 48104 1551 48106
rect 0 48048 1490 48104
rect 1546 48048 1551 48104
rect 0 48046 1551 48048
rect 0 48016 800 48046
rect 1485 48043 1551 48046
rect 4207 47904 4527 47905
rect 4207 47840 4215 47904
rect 4279 47840 4295 47904
rect 4359 47840 4375 47904
rect 4439 47840 4455 47904
rect 4519 47840 4527 47904
rect 4207 47839 4527 47840
rect 7471 47904 7791 47905
rect 7471 47840 7479 47904
rect 7543 47840 7559 47904
rect 7623 47840 7639 47904
rect 7703 47840 7719 47904
rect 7783 47840 7791 47904
rect 7471 47839 7791 47840
rect 10133 47834 10199 47837
rect 11200 47834 12000 47864
rect 10133 47832 12000 47834
rect 10133 47776 10138 47832
rect 10194 47776 12000 47832
rect 10133 47774 12000 47776
rect 10133 47771 10199 47774
rect 11200 47744 12000 47774
rect 0 47562 800 47592
rect 1485 47562 1551 47565
rect 0 47560 1551 47562
rect 0 47504 1490 47560
rect 1546 47504 1551 47560
rect 0 47502 1551 47504
rect 0 47472 800 47502
rect 1485 47499 1551 47502
rect 2576 47360 2896 47361
rect 2576 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2576 47295 2896 47296
rect 5839 47360 6159 47361
rect 5839 47296 5847 47360
rect 5911 47296 5927 47360
rect 5991 47296 6007 47360
rect 6071 47296 6087 47360
rect 6151 47296 6159 47360
rect 5839 47295 6159 47296
rect 9103 47360 9423 47361
rect 9103 47296 9111 47360
rect 9175 47296 9191 47360
rect 9255 47296 9271 47360
rect 9335 47296 9351 47360
rect 9415 47296 9423 47360
rect 9103 47295 9423 47296
rect 3969 47156 4035 47157
rect 3918 47092 3924 47156
rect 3988 47154 4035 47156
rect 3988 47152 4080 47154
rect 4030 47096 4080 47152
rect 3988 47094 4080 47096
rect 3988 47092 4035 47094
rect 3969 47091 4035 47092
rect 0 47018 800 47048
rect 1485 47018 1551 47021
rect 0 47016 1551 47018
rect 0 46960 1490 47016
rect 1546 46960 1551 47016
rect 0 46958 1551 46960
rect 0 46928 800 46958
rect 1485 46955 1551 46958
rect 10133 47018 10199 47021
rect 11200 47018 12000 47048
rect 10133 47016 12000 47018
rect 10133 46960 10138 47016
rect 10194 46960 12000 47016
rect 10133 46958 12000 46960
rect 10133 46955 10199 46958
rect 11200 46928 12000 46958
rect 4207 46816 4527 46817
rect 4207 46752 4215 46816
rect 4279 46752 4295 46816
rect 4359 46752 4375 46816
rect 4439 46752 4455 46816
rect 4519 46752 4527 46816
rect 4207 46751 4527 46752
rect 7471 46816 7791 46817
rect 7471 46752 7479 46816
rect 7543 46752 7559 46816
rect 7623 46752 7639 46816
rect 7703 46752 7719 46816
rect 7783 46752 7791 46816
rect 7471 46751 7791 46752
rect 0 46338 800 46368
rect 1485 46338 1551 46341
rect 3601 46338 3667 46341
rect 0 46336 1551 46338
rect 0 46280 1490 46336
rect 1546 46280 1551 46336
rect 0 46278 1551 46280
rect 0 46248 800 46278
rect 1485 46275 1551 46278
rect 3006 46336 3667 46338
rect 3006 46280 3606 46336
rect 3662 46280 3667 46336
rect 3006 46278 3667 46280
rect 2576 46272 2896 46273
rect 2576 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2576 46207 2896 46208
rect 2681 46066 2747 46069
rect 3006 46066 3066 46278
rect 3601 46275 3667 46278
rect 10133 46338 10199 46341
rect 11200 46338 12000 46368
rect 10133 46336 12000 46338
rect 10133 46280 10138 46336
rect 10194 46280 12000 46336
rect 10133 46278 12000 46280
rect 10133 46275 10199 46278
rect 5839 46272 6159 46273
rect 5839 46208 5847 46272
rect 5911 46208 5927 46272
rect 5991 46208 6007 46272
rect 6071 46208 6087 46272
rect 6151 46208 6159 46272
rect 5839 46207 6159 46208
rect 9103 46272 9423 46273
rect 9103 46208 9111 46272
rect 9175 46208 9191 46272
rect 9255 46208 9271 46272
rect 9335 46208 9351 46272
rect 9415 46208 9423 46272
rect 11200 46248 12000 46278
rect 9103 46207 9423 46208
rect 2681 46064 3066 46066
rect 2681 46008 2686 46064
rect 2742 46008 3066 46064
rect 2681 46006 3066 46008
rect 2681 46003 2747 46006
rect 0 45794 800 45824
rect 1485 45794 1551 45797
rect 0 45792 1551 45794
rect 0 45736 1490 45792
rect 1546 45736 1551 45792
rect 0 45734 1551 45736
rect 0 45704 800 45734
rect 1485 45731 1551 45734
rect 4207 45728 4527 45729
rect 4207 45664 4215 45728
rect 4279 45664 4295 45728
rect 4359 45664 4375 45728
rect 4439 45664 4455 45728
rect 4519 45664 4527 45728
rect 4207 45663 4527 45664
rect 7471 45728 7791 45729
rect 7471 45664 7479 45728
rect 7543 45664 7559 45728
rect 7623 45664 7639 45728
rect 7703 45664 7719 45728
rect 7783 45664 7791 45728
rect 7471 45663 7791 45664
rect 3233 45522 3299 45525
rect 3190 45520 3299 45522
rect 3190 45464 3238 45520
rect 3294 45464 3299 45520
rect 3190 45459 3299 45464
rect 10133 45522 10199 45525
rect 11200 45522 12000 45552
rect 10133 45520 12000 45522
rect 10133 45464 10138 45520
rect 10194 45464 12000 45520
rect 10133 45462 12000 45464
rect 10133 45459 10199 45462
rect 0 45250 800 45280
rect 1485 45250 1551 45253
rect 0 45248 1551 45250
rect 0 45192 1490 45248
rect 1546 45192 1551 45248
rect 0 45190 1551 45192
rect 0 45160 800 45190
rect 1485 45187 1551 45190
rect 2576 45184 2896 45185
rect 2576 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2576 45119 2896 45120
rect 3190 45117 3250 45459
rect 11200 45432 12000 45462
rect 5839 45184 6159 45185
rect 5839 45120 5847 45184
rect 5911 45120 5927 45184
rect 5991 45120 6007 45184
rect 6071 45120 6087 45184
rect 6151 45120 6159 45184
rect 5839 45119 6159 45120
rect 9103 45184 9423 45185
rect 9103 45120 9111 45184
rect 9175 45120 9191 45184
rect 9255 45120 9271 45184
rect 9335 45120 9351 45184
rect 9415 45120 9423 45184
rect 9103 45119 9423 45120
rect 3190 45112 3299 45117
rect 3969 45116 4035 45117
rect 3918 45114 3924 45116
rect 3190 45056 3238 45112
rect 3294 45056 3299 45112
rect 3190 45054 3299 45056
rect 3878 45054 3924 45114
rect 3988 45112 4035 45116
rect 4030 45056 4035 45112
rect 3233 45051 3299 45054
rect 3918 45052 3924 45054
rect 3988 45052 4035 45056
rect 3969 45051 4035 45052
rect 10133 44842 10199 44845
rect 11200 44842 12000 44872
rect 10133 44840 12000 44842
rect 10133 44784 10138 44840
rect 10194 44784 12000 44840
rect 10133 44782 12000 44784
rect 10133 44779 10199 44782
rect 11200 44752 12000 44782
rect 0 44706 800 44736
rect 1485 44706 1551 44709
rect 0 44704 1551 44706
rect 0 44648 1490 44704
rect 1546 44648 1551 44704
rect 0 44646 1551 44648
rect 0 44616 800 44646
rect 1485 44643 1551 44646
rect 4207 44640 4527 44641
rect 4207 44576 4215 44640
rect 4279 44576 4295 44640
rect 4359 44576 4375 44640
rect 4439 44576 4455 44640
rect 4519 44576 4527 44640
rect 4207 44575 4527 44576
rect 7471 44640 7791 44641
rect 7471 44576 7479 44640
rect 7543 44576 7559 44640
rect 7623 44576 7639 44640
rect 7703 44576 7719 44640
rect 7783 44576 7791 44640
rect 7471 44575 7791 44576
rect 0 44162 800 44192
rect 1485 44162 1551 44165
rect 0 44160 1551 44162
rect 0 44104 1490 44160
rect 1546 44104 1551 44160
rect 0 44102 1551 44104
rect 0 44072 800 44102
rect 1485 44099 1551 44102
rect 2576 44096 2896 44097
rect 2576 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2576 44031 2896 44032
rect 5839 44096 6159 44097
rect 5839 44032 5847 44096
rect 5911 44032 5927 44096
rect 5991 44032 6007 44096
rect 6071 44032 6087 44096
rect 6151 44032 6159 44096
rect 5839 44031 6159 44032
rect 9103 44096 9423 44097
rect 9103 44032 9111 44096
rect 9175 44032 9191 44096
rect 9255 44032 9271 44096
rect 9335 44032 9351 44096
rect 9415 44032 9423 44096
rect 9103 44031 9423 44032
rect 10133 44026 10199 44029
rect 11200 44026 12000 44056
rect 10133 44024 12000 44026
rect 10133 43968 10138 44024
rect 10194 43968 12000 44024
rect 10133 43966 12000 43968
rect 10133 43963 10199 43966
rect 11200 43936 12000 43966
rect 0 43618 800 43648
rect 1485 43618 1551 43621
rect 0 43616 1551 43618
rect 0 43560 1490 43616
rect 1546 43560 1551 43616
rect 0 43558 1551 43560
rect 0 43528 800 43558
rect 1485 43555 1551 43558
rect 4207 43552 4527 43553
rect 4207 43488 4215 43552
rect 4279 43488 4295 43552
rect 4359 43488 4375 43552
rect 4439 43488 4455 43552
rect 4519 43488 4527 43552
rect 4207 43487 4527 43488
rect 7471 43552 7791 43553
rect 7471 43488 7479 43552
rect 7543 43488 7559 43552
rect 7623 43488 7639 43552
rect 7703 43488 7719 43552
rect 7783 43488 7791 43552
rect 7471 43487 7791 43488
rect 10133 43346 10199 43349
rect 11200 43346 12000 43376
rect 10133 43344 12000 43346
rect 10133 43288 10138 43344
rect 10194 43288 12000 43344
rect 10133 43286 12000 43288
rect 10133 43283 10199 43286
rect 11200 43256 12000 43286
rect 0 43074 800 43104
rect 1485 43074 1551 43077
rect 0 43072 1551 43074
rect 0 43016 1490 43072
rect 1546 43016 1551 43072
rect 0 43014 1551 43016
rect 0 42984 800 43014
rect 1485 43011 1551 43014
rect 2576 43008 2896 43009
rect 2576 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2576 42943 2896 42944
rect 5839 43008 6159 43009
rect 5839 42944 5847 43008
rect 5911 42944 5927 43008
rect 5991 42944 6007 43008
rect 6071 42944 6087 43008
rect 6151 42944 6159 43008
rect 5839 42943 6159 42944
rect 9103 43008 9423 43009
rect 9103 42944 9111 43008
rect 9175 42944 9191 43008
rect 9255 42944 9271 43008
rect 9335 42944 9351 43008
rect 9415 42944 9423 43008
rect 9103 42943 9423 42944
rect 0 42530 800 42560
rect 1485 42530 1551 42533
rect 0 42528 1551 42530
rect 0 42472 1490 42528
rect 1546 42472 1551 42528
rect 0 42470 1551 42472
rect 0 42440 800 42470
rect 1485 42467 1551 42470
rect 10133 42530 10199 42533
rect 11200 42530 12000 42560
rect 10133 42528 12000 42530
rect 10133 42472 10138 42528
rect 10194 42472 12000 42528
rect 10133 42470 12000 42472
rect 10133 42467 10199 42470
rect 4207 42464 4527 42465
rect 4207 42400 4215 42464
rect 4279 42400 4295 42464
rect 4359 42400 4375 42464
rect 4439 42400 4455 42464
rect 4519 42400 4527 42464
rect 4207 42399 4527 42400
rect 7471 42464 7791 42465
rect 7471 42400 7479 42464
rect 7543 42400 7559 42464
rect 7623 42400 7639 42464
rect 7703 42400 7719 42464
rect 7783 42400 7791 42464
rect 11200 42440 12000 42470
rect 7471 42399 7791 42400
rect 0 41986 800 42016
rect 1485 41986 1551 41989
rect 0 41984 1551 41986
rect 0 41928 1490 41984
rect 1546 41928 1551 41984
rect 0 41926 1551 41928
rect 0 41896 800 41926
rect 1485 41923 1551 41926
rect 2576 41920 2896 41921
rect 2576 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2576 41855 2896 41856
rect 5839 41920 6159 41921
rect 5839 41856 5847 41920
rect 5911 41856 5927 41920
rect 5991 41856 6007 41920
rect 6071 41856 6087 41920
rect 6151 41856 6159 41920
rect 5839 41855 6159 41856
rect 9103 41920 9423 41921
rect 9103 41856 9111 41920
rect 9175 41856 9191 41920
rect 9255 41856 9271 41920
rect 9335 41856 9351 41920
rect 9415 41856 9423 41920
rect 9103 41855 9423 41856
rect 2998 41788 3004 41852
rect 3068 41850 3074 41852
rect 4061 41850 4127 41853
rect 3068 41848 4127 41850
rect 3068 41792 4066 41848
rect 4122 41792 4127 41848
rect 3068 41790 4127 41792
rect 3068 41788 3074 41790
rect 4061 41787 4127 41790
rect 10133 41850 10199 41853
rect 11200 41850 12000 41880
rect 10133 41848 12000 41850
rect 10133 41792 10138 41848
rect 10194 41792 12000 41848
rect 10133 41790 12000 41792
rect 10133 41787 10199 41790
rect 11200 41760 12000 41790
rect 2129 41714 2195 41717
rect 2129 41712 2560 41714
rect 2129 41656 2134 41712
rect 2190 41656 2560 41712
rect 2129 41654 2560 41656
rect 2129 41651 2195 41654
rect 2500 41581 2560 41654
rect 2497 41576 2563 41581
rect 2497 41520 2502 41576
rect 2558 41520 2563 41576
rect 2497 41515 2563 41520
rect 4153 41578 4219 41581
rect 4654 41578 4660 41580
rect 4153 41576 4660 41578
rect 4153 41520 4158 41576
rect 4214 41520 4660 41576
rect 4153 41518 4660 41520
rect 4153 41515 4219 41518
rect 4654 41516 4660 41518
rect 4724 41516 4730 41580
rect 0 41442 800 41472
rect 1485 41442 1551 41445
rect 0 41440 1551 41442
rect 0 41384 1490 41440
rect 1546 41384 1551 41440
rect 0 41382 1551 41384
rect 0 41352 800 41382
rect 1485 41379 1551 41382
rect 4207 41376 4527 41377
rect 4207 41312 4215 41376
rect 4279 41312 4295 41376
rect 4359 41312 4375 41376
rect 4439 41312 4455 41376
rect 4519 41312 4527 41376
rect 4207 41311 4527 41312
rect 7471 41376 7791 41377
rect 7471 41312 7479 41376
rect 7543 41312 7559 41376
rect 7623 41312 7639 41376
rect 7703 41312 7719 41376
rect 7783 41312 7791 41376
rect 7471 41311 7791 41312
rect 2313 41306 2379 41309
rect 2086 41304 2379 41306
rect 2086 41248 2318 41304
rect 2374 41248 2379 41304
rect 2086 41246 2379 41248
rect 1945 41170 2011 41173
rect 2086 41170 2146 41246
rect 2313 41243 2379 41246
rect 6494 41244 6500 41308
rect 6564 41306 6570 41308
rect 6637 41306 6703 41309
rect 6564 41304 6703 41306
rect 6564 41248 6642 41304
rect 6698 41248 6703 41304
rect 6564 41246 6703 41248
rect 6564 41244 6570 41246
rect 6637 41243 6703 41246
rect 1945 41168 2146 41170
rect 1945 41112 1950 41168
rect 2006 41112 2146 41168
rect 1945 41110 2146 41112
rect 2313 41170 2379 41173
rect 2497 41170 2563 41173
rect 2313 41168 2563 41170
rect 2313 41112 2318 41168
rect 2374 41112 2502 41168
rect 2558 41112 2563 41168
rect 2313 41110 2563 41112
rect 1945 41107 2011 41110
rect 2313 41107 2379 41110
rect 2497 41107 2563 41110
rect 2773 41170 2839 41173
rect 4521 41170 4587 41173
rect 2773 41168 4587 41170
rect 2773 41112 2778 41168
rect 2834 41112 4526 41168
rect 4582 41112 4587 41168
rect 2773 41110 4587 41112
rect 2773 41107 2839 41110
rect 4521 41107 4587 41110
rect 10133 41034 10199 41037
rect 11200 41034 12000 41064
rect 10133 41032 12000 41034
rect 10133 40976 10138 41032
rect 10194 40976 12000 41032
rect 10133 40974 12000 40976
rect 10133 40971 10199 40974
rect 11200 40944 12000 40974
rect 0 40898 800 40928
rect 1485 40898 1551 40901
rect 0 40896 1551 40898
rect 0 40840 1490 40896
rect 1546 40840 1551 40896
rect 0 40838 1551 40840
rect 0 40808 800 40838
rect 1485 40835 1551 40838
rect 2576 40832 2896 40833
rect 2576 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2576 40767 2896 40768
rect 5839 40832 6159 40833
rect 5839 40768 5847 40832
rect 5911 40768 5927 40832
rect 5991 40768 6007 40832
rect 6071 40768 6087 40832
rect 6151 40768 6159 40832
rect 5839 40767 6159 40768
rect 9103 40832 9423 40833
rect 9103 40768 9111 40832
rect 9175 40768 9191 40832
rect 9255 40768 9271 40832
rect 9335 40768 9351 40832
rect 9415 40768 9423 40832
rect 9103 40767 9423 40768
rect 0 40354 800 40384
rect 1485 40354 1551 40357
rect 0 40352 1551 40354
rect 0 40296 1490 40352
rect 1546 40296 1551 40352
rect 0 40294 1551 40296
rect 0 40264 800 40294
rect 1485 40291 1551 40294
rect 10133 40354 10199 40357
rect 11200 40354 12000 40384
rect 10133 40352 12000 40354
rect 10133 40296 10138 40352
rect 10194 40296 12000 40352
rect 10133 40294 12000 40296
rect 10133 40291 10199 40294
rect 4207 40288 4527 40289
rect 4207 40224 4215 40288
rect 4279 40224 4295 40288
rect 4359 40224 4375 40288
rect 4439 40224 4455 40288
rect 4519 40224 4527 40288
rect 4207 40223 4527 40224
rect 7471 40288 7791 40289
rect 7471 40224 7479 40288
rect 7543 40224 7559 40288
rect 7623 40224 7639 40288
rect 7703 40224 7719 40288
rect 7783 40224 7791 40288
rect 11200 40264 12000 40294
rect 7471 40223 7791 40224
rect 2589 40082 2655 40085
rect 3049 40084 3115 40085
rect 2998 40082 3004 40084
rect 2589 40080 3004 40082
rect 3068 40082 3115 40084
rect 3068 40080 3196 40082
rect 2589 40024 2594 40080
rect 2650 40024 3004 40080
rect 3110 40024 3196 40080
rect 2589 40022 3004 40024
rect 2589 40019 2655 40022
rect 2998 40020 3004 40022
rect 3068 40022 3196 40024
rect 3068 40020 3115 40022
rect 3049 40019 3115 40020
rect 5073 39946 5139 39949
rect 5073 39944 5274 39946
rect 5073 39888 5078 39944
rect 5134 39888 5274 39944
rect 5073 39886 5274 39888
rect 5073 39883 5139 39886
rect 2576 39744 2896 39745
rect 0 39674 800 39704
rect 2576 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2576 39679 2896 39680
rect 1393 39674 1459 39677
rect 0 39672 1459 39674
rect 0 39616 1398 39672
rect 1454 39616 1459 39672
rect 0 39614 1459 39616
rect 0 39584 800 39614
rect 1393 39611 1459 39614
rect 5214 39405 5274 39886
rect 5839 39744 6159 39745
rect 5839 39680 5847 39744
rect 5911 39680 5927 39744
rect 5991 39680 6007 39744
rect 6071 39680 6087 39744
rect 6151 39680 6159 39744
rect 5839 39679 6159 39680
rect 9103 39744 9423 39745
rect 9103 39680 9111 39744
rect 9175 39680 9191 39744
rect 9255 39680 9271 39744
rect 9335 39680 9351 39744
rect 9415 39680 9423 39744
rect 9103 39679 9423 39680
rect 10133 39538 10199 39541
rect 11200 39538 12000 39568
rect 10133 39536 12000 39538
rect 10133 39480 10138 39536
rect 10194 39480 12000 39536
rect 10133 39478 12000 39480
rect 10133 39475 10199 39478
rect 11200 39448 12000 39478
rect 5214 39400 5323 39405
rect 5214 39344 5262 39400
rect 5318 39344 5323 39400
rect 5214 39342 5323 39344
rect 5257 39339 5323 39342
rect 4207 39200 4527 39201
rect 0 39130 800 39160
rect 4207 39136 4215 39200
rect 4279 39136 4295 39200
rect 4359 39136 4375 39200
rect 4439 39136 4455 39200
rect 4519 39136 4527 39200
rect 4207 39135 4527 39136
rect 7471 39200 7791 39201
rect 7471 39136 7479 39200
rect 7543 39136 7559 39200
rect 7623 39136 7639 39200
rect 7703 39136 7719 39200
rect 7783 39136 7791 39200
rect 7471 39135 7791 39136
rect 1393 39130 1459 39133
rect 0 39128 1459 39130
rect 0 39072 1398 39128
rect 1454 39072 1459 39128
rect 0 39070 1459 39072
rect 0 39040 800 39070
rect 1393 39067 1459 39070
rect 10133 38722 10199 38725
rect 11200 38722 12000 38752
rect 10133 38720 12000 38722
rect 10133 38664 10138 38720
rect 10194 38664 12000 38720
rect 10133 38662 12000 38664
rect 10133 38659 10199 38662
rect 2576 38656 2896 38657
rect 0 38586 800 38616
rect 2576 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2576 38591 2896 38592
rect 5839 38656 6159 38657
rect 5839 38592 5847 38656
rect 5911 38592 5927 38656
rect 5991 38592 6007 38656
rect 6071 38592 6087 38656
rect 6151 38592 6159 38656
rect 5839 38591 6159 38592
rect 9103 38656 9423 38657
rect 9103 38592 9111 38656
rect 9175 38592 9191 38656
rect 9255 38592 9271 38656
rect 9335 38592 9351 38656
rect 9415 38592 9423 38656
rect 11200 38632 12000 38662
rect 9103 38591 9423 38592
rect 1393 38586 1459 38589
rect 0 38584 1459 38586
rect 0 38528 1398 38584
rect 1454 38528 1459 38584
rect 0 38526 1459 38528
rect 0 38496 800 38526
rect 1393 38523 1459 38526
rect 4207 38112 4527 38113
rect 0 38042 800 38072
rect 4207 38048 4215 38112
rect 4279 38048 4295 38112
rect 4359 38048 4375 38112
rect 4439 38048 4455 38112
rect 4519 38048 4527 38112
rect 4207 38047 4527 38048
rect 7471 38112 7791 38113
rect 7471 38048 7479 38112
rect 7543 38048 7559 38112
rect 7623 38048 7639 38112
rect 7703 38048 7719 38112
rect 7783 38048 7791 38112
rect 7471 38047 7791 38048
rect 1393 38042 1459 38045
rect 0 38040 1459 38042
rect 0 37984 1398 38040
rect 1454 37984 1459 38040
rect 0 37982 1459 37984
rect 0 37952 800 37982
rect 1393 37979 1459 37982
rect 10133 38042 10199 38045
rect 11200 38042 12000 38072
rect 10133 38040 12000 38042
rect 10133 37984 10138 38040
rect 10194 37984 12000 38040
rect 10133 37982 12000 37984
rect 10133 37979 10199 37982
rect 11200 37952 12000 37982
rect 2576 37568 2896 37569
rect 0 37498 800 37528
rect 2576 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2576 37503 2896 37504
rect 5839 37568 6159 37569
rect 5839 37504 5847 37568
rect 5911 37504 5927 37568
rect 5991 37504 6007 37568
rect 6071 37504 6087 37568
rect 6151 37504 6159 37568
rect 5839 37503 6159 37504
rect 9103 37568 9423 37569
rect 9103 37504 9111 37568
rect 9175 37504 9191 37568
rect 9255 37504 9271 37568
rect 9335 37504 9351 37568
rect 9415 37504 9423 37568
rect 9103 37503 9423 37504
rect 1393 37498 1459 37501
rect 0 37496 1459 37498
rect 0 37440 1398 37496
rect 1454 37440 1459 37496
rect 0 37438 1459 37440
rect 0 37408 800 37438
rect 1393 37435 1459 37438
rect 10133 37226 10199 37229
rect 11200 37226 12000 37256
rect 10133 37224 12000 37226
rect 10133 37168 10138 37224
rect 10194 37168 12000 37224
rect 10133 37166 12000 37168
rect 10133 37163 10199 37166
rect 11200 37136 12000 37166
rect 4207 37024 4527 37025
rect 0 36954 800 36984
rect 4207 36960 4215 37024
rect 4279 36960 4295 37024
rect 4359 36960 4375 37024
rect 4439 36960 4455 37024
rect 4519 36960 4527 37024
rect 4207 36959 4527 36960
rect 7471 37024 7791 37025
rect 7471 36960 7479 37024
rect 7543 36960 7559 37024
rect 7623 36960 7639 37024
rect 7703 36960 7719 37024
rect 7783 36960 7791 37024
rect 7471 36959 7791 36960
rect 1393 36954 1459 36957
rect 6453 36956 6519 36957
rect 6453 36954 6500 36956
rect 0 36952 1459 36954
rect 0 36896 1398 36952
rect 1454 36896 1459 36952
rect 0 36894 1459 36896
rect 6408 36952 6500 36954
rect 6408 36896 6458 36952
rect 6408 36894 6500 36896
rect 0 36864 800 36894
rect 1393 36891 1459 36894
rect 6453 36892 6500 36894
rect 6564 36892 6570 36956
rect 6453 36891 6519 36892
rect 10133 36546 10199 36549
rect 11200 36546 12000 36576
rect 10133 36544 12000 36546
rect 10133 36488 10138 36544
rect 10194 36488 12000 36544
rect 10133 36486 12000 36488
rect 10133 36483 10199 36486
rect 2576 36480 2896 36481
rect 0 36410 800 36440
rect 2576 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2576 36415 2896 36416
rect 5839 36480 6159 36481
rect 5839 36416 5847 36480
rect 5911 36416 5927 36480
rect 5991 36416 6007 36480
rect 6071 36416 6087 36480
rect 6151 36416 6159 36480
rect 5839 36415 6159 36416
rect 9103 36480 9423 36481
rect 9103 36416 9111 36480
rect 9175 36416 9191 36480
rect 9255 36416 9271 36480
rect 9335 36416 9351 36480
rect 9415 36416 9423 36480
rect 11200 36456 12000 36486
rect 9103 36415 9423 36416
rect 1393 36410 1459 36413
rect 0 36408 1459 36410
rect 0 36352 1398 36408
rect 1454 36352 1459 36408
rect 0 36350 1459 36352
rect 0 36320 800 36350
rect 1393 36347 1459 36350
rect 4207 35936 4527 35937
rect 0 35866 800 35896
rect 4207 35872 4215 35936
rect 4279 35872 4295 35936
rect 4359 35872 4375 35936
rect 4439 35872 4455 35936
rect 4519 35872 4527 35936
rect 4207 35871 4527 35872
rect 7471 35936 7791 35937
rect 7471 35872 7479 35936
rect 7543 35872 7559 35936
rect 7623 35872 7639 35936
rect 7703 35872 7719 35936
rect 7783 35872 7791 35936
rect 7471 35871 7791 35872
rect 1393 35866 1459 35869
rect 5349 35866 5415 35869
rect 0 35864 1459 35866
rect 0 35808 1398 35864
rect 1454 35808 1459 35864
rect 0 35806 1459 35808
rect 0 35776 800 35806
rect 1393 35803 1459 35806
rect 5214 35864 5415 35866
rect 5214 35808 5354 35864
rect 5410 35808 5415 35864
rect 5214 35806 5415 35808
rect 5073 35458 5139 35461
rect 5214 35458 5274 35806
rect 5349 35803 5415 35806
rect 10133 35730 10199 35733
rect 11200 35730 12000 35760
rect 10133 35728 12000 35730
rect 10133 35672 10138 35728
rect 10194 35672 12000 35728
rect 10133 35670 12000 35672
rect 10133 35667 10199 35670
rect 11200 35640 12000 35670
rect 5073 35456 5274 35458
rect 5073 35400 5078 35456
rect 5134 35400 5274 35456
rect 5073 35398 5274 35400
rect 5073 35395 5139 35398
rect 2576 35392 2896 35393
rect 0 35322 800 35352
rect 2576 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2576 35327 2896 35328
rect 5839 35392 6159 35393
rect 5839 35328 5847 35392
rect 5911 35328 5927 35392
rect 5991 35328 6007 35392
rect 6071 35328 6087 35392
rect 6151 35328 6159 35392
rect 5839 35327 6159 35328
rect 9103 35392 9423 35393
rect 9103 35328 9111 35392
rect 9175 35328 9191 35392
rect 9255 35328 9271 35392
rect 9335 35328 9351 35392
rect 9415 35328 9423 35392
rect 9103 35327 9423 35328
rect 1393 35322 1459 35325
rect 0 35320 1459 35322
rect 0 35264 1398 35320
rect 1454 35264 1459 35320
rect 0 35262 1459 35264
rect 0 35232 800 35262
rect 1393 35259 1459 35262
rect 10133 35050 10199 35053
rect 11200 35050 12000 35080
rect 10133 35048 12000 35050
rect 10133 34992 10138 35048
rect 10194 34992 12000 35048
rect 10133 34990 12000 34992
rect 10133 34987 10199 34990
rect 11200 34960 12000 34990
rect 4207 34848 4527 34849
rect 0 34778 800 34808
rect 4207 34784 4215 34848
rect 4279 34784 4295 34848
rect 4359 34784 4375 34848
rect 4439 34784 4455 34848
rect 4519 34784 4527 34848
rect 4207 34783 4527 34784
rect 7471 34848 7791 34849
rect 7471 34784 7479 34848
rect 7543 34784 7559 34848
rect 7623 34784 7639 34848
rect 7703 34784 7719 34848
rect 7783 34784 7791 34848
rect 7471 34783 7791 34784
rect 1393 34778 1459 34781
rect 0 34776 1459 34778
rect 0 34720 1398 34776
rect 1454 34720 1459 34776
rect 0 34718 1459 34720
rect 0 34688 800 34718
rect 1393 34715 1459 34718
rect 4613 34372 4679 34373
rect 4613 34368 4660 34372
rect 4724 34370 4730 34372
rect 4613 34312 4618 34368
rect 4613 34308 4660 34312
rect 4724 34310 4770 34370
rect 4724 34308 4730 34310
rect 4613 34307 4679 34308
rect 2576 34304 2896 34305
rect 0 34234 800 34264
rect 2576 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2576 34239 2896 34240
rect 5839 34304 6159 34305
rect 5839 34240 5847 34304
rect 5911 34240 5927 34304
rect 5991 34240 6007 34304
rect 6071 34240 6087 34304
rect 6151 34240 6159 34304
rect 5839 34239 6159 34240
rect 9103 34304 9423 34305
rect 9103 34240 9111 34304
rect 9175 34240 9191 34304
rect 9255 34240 9271 34304
rect 9335 34240 9351 34304
rect 9415 34240 9423 34304
rect 9103 34239 9423 34240
rect 1393 34234 1459 34237
rect 0 34232 1459 34234
rect 0 34176 1398 34232
rect 1454 34176 1459 34232
rect 0 34174 1459 34176
rect 0 34144 800 34174
rect 1393 34171 1459 34174
rect 10133 34234 10199 34237
rect 11200 34234 12000 34264
rect 10133 34232 12000 34234
rect 10133 34176 10138 34232
rect 10194 34176 12000 34232
rect 10133 34174 12000 34176
rect 10133 34171 10199 34174
rect 11200 34144 12000 34174
rect 4207 33760 4527 33761
rect 0 33690 800 33720
rect 4207 33696 4215 33760
rect 4279 33696 4295 33760
rect 4359 33696 4375 33760
rect 4439 33696 4455 33760
rect 4519 33696 4527 33760
rect 4207 33695 4527 33696
rect 7471 33760 7791 33761
rect 7471 33696 7479 33760
rect 7543 33696 7559 33760
rect 7623 33696 7639 33760
rect 7703 33696 7719 33760
rect 7783 33696 7791 33760
rect 7471 33695 7791 33696
rect 1393 33690 1459 33693
rect 0 33688 1459 33690
rect 0 33632 1398 33688
rect 1454 33632 1459 33688
rect 0 33630 1459 33632
rect 0 33600 800 33630
rect 1393 33627 1459 33630
rect 10133 33554 10199 33557
rect 11200 33554 12000 33584
rect 10133 33552 12000 33554
rect 10133 33496 10138 33552
rect 10194 33496 12000 33552
rect 10133 33494 12000 33496
rect 10133 33491 10199 33494
rect 11200 33464 12000 33494
rect 2576 33216 2896 33217
rect 2576 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2576 33151 2896 33152
rect 5839 33216 6159 33217
rect 5839 33152 5847 33216
rect 5911 33152 5927 33216
rect 5991 33152 6007 33216
rect 6071 33152 6087 33216
rect 6151 33152 6159 33216
rect 5839 33151 6159 33152
rect 9103 33216 9423 33217
rect 9103 33152 9111 33216
rect 9175 33152 9191 33216
rect 9255 33152 9271 33216
rect 9335 33152 9351 33216
rect 9415 33152 9423 33216
rect 9103 33151 9423 33152
rect 0 33010 800 33040
rect 1393 33010 1459 33013
rect 0 33008 1459 33010
rect 0 32952 1398 33008
rect 1454 32952 1459 33008
rect 0 32950 1459 32952
rect 0 32920 800 32950
rect 1393 32947 1459 32950
rect 10133 32738 10199 32741
rect 11200 32738 12000 32768
rect 10133 32736 12000 32738
rect 10133 32680 10138 32736
rect 10194 32680 12000 32736
rect 10133 32678 12000 32680
rect 10133 32675 10199 32678
rect 4207 32672 4527 32673
rect 4207 32608 4215 32672
rect 4279 32608 4295 32672
rect 4359 32608 4375 32672
rect 4439 32608 4455 32672
rect 4519 32608 4527 32672
rect 4207 32607 4527 32608
rect 7471 32672 7791 32673
rect 7471 32608 7479 32672
rect 7543 32608 7559 32672
rect 7623 32608 7639 32672
rect 7703 32608 7719 32672
rect 7783 32608 7791 32672
rect 11200 32648 12000 32678
rect 7471 32607 7791 32608
rect 0 32466 800 32496
rect 1393 32466 1459 32469
rect 0 32464 1459 32466
rect 0 32408 1398 32464
rect 1454 32408 1459 32464
rect 0 32406 1459 32408
rect 0 32376 800 32406
rect 1393 32403 1459 32406
rect 2576 32128 2896 32129
rect 2576 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2576 32063 2896 32064
rect 5839 32128 6159 32129
rect 5839 32064 5847 32128
rect 5911 32064 5927 32128
rect 5991 32064 6007 32128
rect 6071 32064 6087 32128
rect 6151 32064 6159 32128
rect 5839 32063 6159 32064
rect 9103 32128 9423 32129
rect 9103 32064 9111 32128
rect 9175 32064 9191 32128
rect 9255 32064 9271 32128
rect 9335 32064 9351 32128
rect 9415 32064 9423 32128
rect 9103 32063 9423 32064
rect 0 31922 800 31952
rect 1301 31922 1367 31925
rect 0 31920 1367 31922
rect 0 31864 1306 31920
rect 1362 31864 1367 31920
rect 0 31862 1367 31864
rect 0 31832 800 31862
rect 1301 31859 1367 31862
rect 10133 31922 10199 31925
rect 11200 31922 12000 31952
rect 10133 31920 12000 31922
rect 10133 31864 10138 31920
rect 10194 31864 12000 31920
rect 10133 31862 12000 31864
rect 10133 31859 10199 31862
rect 11200 31832 12000 31862
rect 4207 31584 4527 31585
rect 4207 31520 4215 31584
rect 4279 31520 4295 31584
rect 4359 31520 4375 31584
rect 4439 31520 4455 31584
rect 4519 31520 4527 31584
rect 4207 31519 4527 31520
rect 7471 31584 7791 31585
rect 7471 31520 7479 31584
rect 7543 31520 7559 31584
rect 7623 31520 7639 31584
rect 7703 31520 7719 31584
rect 7783 31520 7791 31584
rect 7471 31519 7791 31520
rect 0 31378 800 31408
rect 1393 31378 1459 31381
rect 0 31376 1459 31378
rect 0 31320 1398 31376
rect 1454 31320 1459 31376
rect 0 31318 1459 31320
rect 0 31288 800 31318
rect 1393 31315 1459 31318
rect 10133 31242 10199 31245
rect 11200 31242 12000 31272
rect 10133 31240 12000 31242
rect 10133 31184 10138 31240
rect 10194 31184 12000 31240
rect 10133 31182 12000 31184
rect 10133 31179 10199 31182
rect 11200 31152 12000 31182
rect 2576 31040 2896 31041
rect 2576 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2576 30975 2896 30976
rect 5839 31040 6159 31041
rect 5839 30976 5847 31040
rect 5911 30976 5927 31040
rect 5991 30976 6007 31040
rect 6071 30976 6087 31040
rect 6151 30976 6159 31040
rect 5839 30975 6159 30976
rect 9103 31040 9423 31041
rect 9103 30976 9111 31040
rect 9175 30976 9191 31040
rect 9255 30976 9271 31040
rect 9335 30976 9351 31040
rect 9415 30976 9423 31040
rect 9103 30975 9423 30976
rect 0 30834 800 30864
rect 1301 30834 1367 30837
rect 0 30832 1367 30834
rect 0 30776 1306 30832
rect 1362 30776 1367 30832
rect 0 30774 1367 30776
rect 0 30744 800 30774
rect 1301 30771 1367 30774
rect 4207 30496 4527 30497
rect 4207 30432 4215 30496
rect 4279 30432 4295 30496
rect 4359 30432 4375 30496
rect 4439 30432 4455 30496
rect 4519 30432 4527 30496
rect 4207 30431 4527 30432
rect 7471 30496 7791 30497
rect 7471 30432 7479 30496
rect 7543 30432 7559 30496
rect 7623 30432 7639 30496
rect 7703 30432 7719 30496
rect 7783 30432 7791 30496
rect 7471 30431 7791 30432
rect 10133 30426 10199 30429
rect 11200 30426 12000 30456
rect 10133 30424 12000 30426
rect 10133 30368 10138 30424
rect 10194 30368 12000 30424
rect 10133 30366 12000 30368
rect 10133 30363 10199 30366
rect 11200 30336 12000 30366
rect 0 30290 800 30320
rect 1393 30290 1459 30293
rect 0 30288 1459 30290
rect 0 30232 1398 30288
rect 1454 30232 1459 30288
rect 0 30230 1459 30232
rect 0 30200 800 30230
rect 1393 30227 1459 30230
rect 2576 29952 2896 29953
rect 2576 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2576 29887 2896 29888
rect 5839 29952 6159 29953
rect 5839 29888 5847 29952
rect 5911 29888 5927 29952
rect 5991 29888 6007 29952
rect 6071 29888 6087 29952
rect 6151 29888 6159 29952
rect 5839 29887 6159 29888
rect 9103 29952 9423 29953
rect 9103 29888 9111 29952
rect 9175 29888 9191 29952
rect 9255 29888 9271 29952
rect 9335 29888 9351 29952
rect 9415 29888 9423 29952
rect 9103 29887 9423 29888
rect 0 29746 800 29776
rect 1301 29746 1367 29749
rect 0 29744 1367 29746
rect 0 29688 1306 29744
rect 1362 29688 1367 29744
rect 0 29686 1367 29688
rect 0 29656 800 29686
rect 1301 29683 1367 29686
rect 10133 29746 10199 29749
rect 11200 29746 12000 29776
rect 10133 29744 12000 29746
rect 10133 29688 10138 29744
rect 10194 29688 12000 29744
rect 10133 29686 12000 29688
rect 10133 29683 10199 29686
rect 11200 29656 12000 29686
rect 4207 29408 4527 29409
rect 4207 29344 4215 29408
rect 4279 29344 4295 29408
rect 4359 29344 4375 29408
rect 4439 29344 4455 29408
rect 4519 29344 4527 29408
rect 4207 29343 4527 29344
rect 7471 29408 7791 29409
rect 7471 29344 7479 29408
rect 7543 29344 7559 29408
rect 7623 29344 7639 29408
rect 7703 29344 7719 29408
rect 7783 29344 7791 29408
rect 7471 29343 7791 29344
rect 0 29202 800 29232
rect 1393 29202 1459 29205
rect 0 29200 1459 29202
rect 0 29144 1398 29200
rect 1454 29144 1459 29200
rect 0 29142 1459 29144
rect 0 29112 800 29142
rect 1393 29139 1459 29142
rect 10133 28930 10199 28933
rect 11200 28930 12000 28960
rect 10133 28928 12000 28930
rect 10133 28872 10138 28928
rect 10194 28872 12000 28928
rect 10133 28870 12000 28872
rect 10133 28867 10199 28870
rect 2576 28864 2896 28865
rect 2576 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2576 28799 2896 28800
rect 5839 28864 6159 28865
rect 5839 28800 5847 28864
rect 5911 28800 5927 28864
rect 5991 28800 6007 28864
rect 6071 28800 6087 28864
rect 6151 28800 6159 28864
rect 5839 28799 6159 28800
rect 9103 28864 9423 28865
rect 9103 28800 9111 28864
rect 9175 28800 9191 28864
rect 9255 28800 9271 28864
rect 9335 28800 9351 28864
rect 9415 28800 9423 28864
rect 11200 28840 12000 28870
rect 9103 28799 9423 28800
rect 0 28658 800 28688
rect 1301 28658 1367 28661
rect 0 28656 1367 28658
rect 0 28600 1306 28656
rect 1362 28600 1367 28656
rect 0 28598 1367 28600
rect 0 28568 800 28598
rect 1301 28595 1367 28598
rect 4207 28320 4527 28321
rect 4207 28256 4215 28320
rect 4279 28256 4295 28320
rect 4359 28256 4375 28320
rect 4439 28256 4455 28320
rect 4519 28256 4527 28320
rect 4207 28255 4527 28256
rect 7471 28320 7791 28321
rect 7471 28256 7479 28320
rect 7543 28256 7559 28320
rect 7623 28256 7639 28320
rect 7703 28256 7719 28320
rect 7783 28256 7791 28320
rect 7471 28255 7791 28256
rect 10133 28250 10199 28253
rect 11200 28250 12000 28280
rect 10133 28248 12000 28250
rect 10133 28192 10138 28248
rect 10194 28192 12000 28248
rect 10133 28190 12000 28192
rect 10133 28187 10199 28190
rect 11200 28160 12000 28190
rect 0 28114 800 28144
rect 1393 28114 1459 28117
rect 0 28112 1459 28114
rect 0 28056 1398 28112
rect 1454 28056 1459 28112
rect 0 28054 1459 28056
rect 0 28024 800 28054
rect 1393 28051 1459 28054
rect 2576 27776 2896 27777
rect 2576 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2576 27711 2896 27712
rect 5839 27776 6159 27777
rect 5839 27712 5847 27776
rect 5911 27712 5927 27776
rect 5991 27712 6007 27776
rect 6071 27712 6087 27776
rect 6151 27712 6159 27776
rect 5839 27711 6159 27712
rect 9103 27776 9423 27777
rect 9103 27712 9111 27776
rect 9175 27712 9191 27776
rect 9255 27712 9271 27776
rect 9335 27712 9351 27776
rect 9415 27712 9423 27776
rect 9103 27711 9423 27712
rect 0 27570 800 27600
rect 1301 27570 1367 27573
rect 0 27568 1367 27570
rect 0 27512 1306 27568
rect 1362 27512 1367 27568
rect 0 27510 1367 27512
rect 0 27480 800 27510
rect 1301 27507 1367 27510
rect 10133 27434 10199 27437
rect 11200 27434 12000 27464
rect 10133 27432 12000 27434
rect 10133 27376 10138 27432
rect 10194 27376 12000 27432
rect 10133 27374 12000 27376
rect 10133 27371 10199 27374
rect 11200 27344 12000 27374
rect 4207 27232 4527 27233
rect 4207 27168 4215 27232
rect 4279 27168 4295 27232
rect 4359 27168 4375 27232
rect 4439 27168 4455 27232
rect 4519 27168 4527 27232
rect 4207 27167 4527 27168
rect 7471 27232 7791 27233
rect 7471 27168 7479 27232
rect 7543 27168 7559 27232
rect 7623 27168 7639 27232
rect 7703 27168 7719 27232
rect 7783 27168 7791 27232
rect 7471 27167 7791 27168
rect 0 27026 800 27056
rect 1945 27026 2011 27029
rect 0 27024 2011 27026
rect 0 26968 1950 27024
rect 2006 26968 2011 27024
rect 0 26966 2011 26968
rect 0 26936 800 26966
rect 1945 26963 2011 26966
rect 10225 26754 10291 26757
rect 11200 26754 12000 26784
rect 10225 26752 12000 26754
rect 10225 26696 10230 26752
rect 10286 26696 12000 26752
rect 10225 26694 12000 26696
rect 10225 26691 10291 26694
rect 2576 26688 2896 26689
rect 2576 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2576 26623 2896 26624
rect 5839 26688 6159 26689
rect 5839 26624 5847 26688
rect 5911 26624 5927 26688
rect 5991 26624 6007 26688
rect 6071 26624 6087 26688
rect 6151 26624 6159 26688
rect 5839 26623 6159 26624
rect 9103 26688 9423 26689
rect 9103 26624 9111 26688
rect 9175 26624 9191 26688
rect 9255 26624 9271 26688
rect 9335 26624 9351 26688
rect 9415 26624 9423 26688
rect 11200 26664 12000 26694
rect 9103 26623 9423 26624
rect 0 26346 800 26376
rect 1945 26346 2011 26349
rect 0 26344 2011 26346
rect 0 26288 1950 26344
rect 2006 26288 2011 26344
rect 0 26286 2011 26288
rect 0 26256 800 26286
rect 1945 26283 2011 26286
rect 4207 26144 4527 26145
rect 4207 26080 4215 26144
rect 4279 26080 4295 26144
rect 4359 26080 4375 26144
rect 4439 26080 4455 26144
rect 4519 26080 4527 26144
rect 4207 26079 4527 26080
rect 7471 26144 7791 26145
rect 7471 26080 7479 26144
rect 7543 26080 7559 26144
rect 7623 26080 7639 26144
rect 7703 26080 7719 26144
rect 7783 26080 7791 26144
rect 7471 26079 7791 26080
rect 10041 25938 10107 25941
rect 11200 25938 12000 25968
rect 10041 25936 12000 25938
rect 10041 25880 10046 25936
rect 10102 25880 12000 25936
rect 10041 25878 12000 25880
rect 10041 25875 10107 25878
rect 11200 25848 12000 25878
rect 0 25802 800 25832
rect 1945 25802 2011 25805
rect 0 25800 2011 25802
rect 0 25744 1950 25800
rect 2006 25744 2011 25800
rect 0 25742 2011 25744
rect 0 25712 800 25742
rect 1945 25739 2011 25742
rect 2576 25600 2896 25601
rect 2576 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2576 25535 2896 25536
rect 5839 25600 6159 25601
rect 5839 25536 5847 25600
rect 5911 25536 5927 25600
rect 5991 25536 6007 25600
rect 6071 25536 6087 25600
rect 6151 25536 6159 25600
rect 5839 25535 6159 25536
rect 9103 25600 9423 25601
rect 9103 25536 9111 25600
rect 9175 25536 9191 25600
rect 9255 25536 9271 25600
rect 9335 25536 9351 25600
rect 9415 25536 9423 25600
rect 9103 25535 9423 25536
rect 0 25258 800 25288
rect 1945 25258 2011 25261
rect 0 25256 2011 25258
rect 0 25200 1950 25256
rect 2006 25200 2011 25256
rect 0 25198 2011 25200
rect 0 25168 800 25198
rect 1945 25195 2011 25198
rect 10133 25258 10199 25261
rect 11200 25258 12000 25288
rect 10133 25256 12000 25258
rect 10133 25200 10138 25256
rect 10194 25200 12000 25256
rect 10133 25198 12000 25200
rect 10133 25195 10199 25198
rect 11200 25168 12000 25198
rect 4207 25056 4527 25057
rect 4207 24992 4215 25056
rect 4279 24992 4295 25056
rect 4359 24992 4375 25056
rect 4439 24992 4455 25056
rect 4519 24992 4527 25056
rect 4207 24991 4527 24992
rect 7471 25056 7791 25057
rect 7471 24992 7479 25056
rect 7543 24992 7559 25056
rect 7623 24992 7639 25056
rect 7703 24992 7719 25056
rect 7783 24992 7791 25056
rect 7471 24991 7791 24992
rect 0 24714 800 24744
rect 1945 24714 2011 24717
rect 0 24712 2011 24714
rect 0 24656 1950 24712
rect 2006 24656 2011 24712
rect 0 24654 2011 24656
rect 0 24624 800 24654
rect 1945 24651 2011 24654
rect 2576 24512 2896 24513
rect 2576 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2576 24447 2896 24448
rect 5839 24512 6159 24513
rect 5839 24448 5847 24512
rect 5911 24448 5927 24512
rect 5991 24448 6007 24512
rect 6071 24448 6087 24512
rect 6151 24448 6159 24512
rect 5839 24447 6159 24448
rect 9103 24512 9423 24513
rect 9103 24448 9111 24512
rect 9175 24448 9191 24512
rect 9255 24448 9271 24512
rect 9335 24448 9351 24512
rect 9415 24448 9423 24512
rect 9103 24447 9423 24448
rect 10133 24442 10199 24445
rect 11200 24442 12000 24472
rect 10133 24440 12000 24442
rect 10133 24384 10138 24440
rect 10194 24384 12000 24440
rect 10133 24382 12000 24384
rect 10133 24379 10199 24382
rect 11200 24352 12000 24382
rect 0 24170 800 24200
rect 1945 24170 2011 24173
rect 0 24168 2011 24170
rect 0 24112 1950 24168
rect 2006 24112 2011 24168
rect 0 24110 2011 24112
rect 0 24080 800 24110
rect 1945 24107 2011 24110
rect 4207 23968 4527 23969
rect 4207 23904 4215 23968
rect 4279 23904 4295 23968
rect 4359 23904 4375 23968
rect 4439 23904 4455 23968
rect 4519 23904 4527 23968
rect 4207 23903 4527 23904
rect 7471 23968 7791 23969
rect 7471 23904 7479 23968
rect 7543 23904 7559 23968
rect 7623 23904 7639 23968
rect 7703 23904 7719 23968
rect 7783 23904 7791 23968
rect 7471 23903 7791 23904
rect 0 23626 800 23656
rect 1853 23626 1919 23629
rect 0 23624 1919 23626
rect 0 23568 1858 23624
rect 1914 23568 1919 23624
rect 0 23566 1919 23568
rect 0 23536 800 23566
rect 1853 23563 1919 23566
rect 10133 23626 10199 23629
rect 11200 23626 12000 23656
rect 10133 23624 12000 23626
rect 10133 23568 10138 23624
rect 10194 23568 12000 23624
rect 10133 23566 12000 23568
rect 10133 23563 10199 23566
rect 11200 23536 12000 23566
rect 2576 23424 2896 23425
rect 2576 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2576 23359 2896 23360
rect 5839 23424 6159 23425
rect 5839 23360 5847 23424
rect 5911 23360 5927 23424
rect 5991 23360 6007 23424
rect 6071 23360 6087 23424
rect 6151 23360 6159 23424
rect 5839 23359 6159 23360
rect 9103 23424 9423 23425
rect 9103 23360 9111 23424
rect 9175 23360 9191 23424
rect 9255 23360 9271 23424
rect 9335 23360 9351 23424
rect 9415 23360 9423 23424
rect 9103 23359 9423 23360
rect 0 23082 800 23112
rect 1945 23082 2011 23085
rect 0 23080 2011 23082
rect 0 23024 1950 23080
rect 2006 23024 2011 23080
rect 0 23022 2011 23024
rect 0 22992 800 23022
rect 1945 23019 2011 23022
rect 9121 22946 9187 22949
rect 11200 22946 12000 22976
rect 9121 22944 12000 22946
rect 9121 22888 9126 22944
rect 9182 22888 12000 22944
rect 9121 22886 12000 22888
rect 9121 22883 9187 22886
rect 4207 22880 4527 22881
rect 4207 22816 4215 22880
rect 4279 22816 4295 22880
rect 4359 22816 4375 22880
rect 4439 22816 4455 22880
rect 4519 22816 4527 22880
rect 4207 22815 4527 22816
rect 7471 22880 7791 22881
rect 7471 22816 7479 22880
rect 7543 22816 7559 22880
rect 7623 22816 7639 22880
rect 7703 22816 7719 22880
rect 7783 22816 7791 22880
rect 11200 22856 12000 22886
rect 7471 22815 7791 22816
rect 0 22538 800 22568
rect 1945 22538 2011 22541
rect 0 22536 2011 22538
rect 0 22480 1950 22536
rect 2006 22480 2011 22536
rect 0 22478 2011 22480
rect 0 22448 800 22478
rect 1945 22475 2011 22478
rect 2576 22336 2896 22337
rect 2576 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2576 22271 2896 22272
rect 5839 22336 6159 22337
rect 5839 22272 5847 22336
rect 5911 22272 5927 22336
rect 5991 22272 6007 22336
rect 6071 22272 6087 22336
rect 6151 22272 6159 22336
rect 5839 22271 6159 22272
rect 9103 22336 9423 22337
rect 9103 22272 9111 22336
rect 9175 22272 9191 22336
rect 9255 22272 9271 22336
rect 9335 22272 9351 22336
rect 9415 22272 9423 22336
rect 9103 22271 9423 22272
rect 8845 22130 8911 22133
rect 11200 22130 12000 22160
rect 8845 22128 12000 22130
rect 8845 22072 8850 22128
rect 8906 22072 12000 22128
rect 8845 22070 12000 22072
rect 8845 22067 8911 22070
rect 11200 22040 12000 22070
rect 0 21994 800 22024
rect 1945 21994 2011 21997
rect 0 21992 2011 21994
rect 0 21936 1950 21992
rect 2006 21936 2011 21992
rect 0 21934 2011 21936
rect 0 21904 800 21934
rect 1945 21931 2011 21934
rect 4207 21792 4527 21793
rect 4207 21728 4215 21792
rect 4279 21728 4295 21792
rect 4359 21728 4375 21792
rect 4439 21728 4455 21792
rect 4519 21728 4527 21792
rect 4207 21727 4527 21728
rect 7471 21792 7791 21793
rect 7471 21728 7479 21792
rect 7543 21728 7559 21792
rect 7623 21728 7639 21792
rect 7703 21728 7719 21792
rect 7783 21728 7791 21792
rect 7471 21727 7791 21728
rect 0 21450 800 21480
rect 1485 21450 1551 21453
rect 0 21448 1551 21450
rect 0 21392 1490 21448
rect 1546 21392 1551 21448
rect 0 21390 1551 21392
rect 0 21360 800 21390
rect 1485 21387 1551 21390
rect 8937 21450 9003 21453
rect 11200 21450 12000 21480
rect 8937 21448 12000 21450
rect 8937 21392 8942 21448
rect 8998 21392 12000 21448
rect 8937 21390 12000 21392
rect 8937 21387 9003 21390
rect 11200 21360 12000 21390
rect 2576 21248 2896 21249
rect 2576 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2576 21183 2896 21184
rect 5839 21248 6159 21249
rect 5839 21184 5847 21248
rect 5911 21184 5927 21248
rect 5991 21184 6007 21248
rect 6071 21184 6087 21248
rect 6151 21184 6159 21248
rect 5839 21183 6159 21184
rect 9103 21248 9423 21249
rect 9103 21184 9111 21248
rect 9175 21184 9191 21248
rect 9255 21184 9271 21248
rect 9335 21184 9351 21248
rect 9415 21184 9423 21248
rect 9103 21183 9423 21184
rect 0 20906 800 20936
rect 1485 20906 1551 20909
rect 0 20904 1551 20906
rect 0 20848 1490 20904
rect 1546 20848 1551 20904
rect 0 20846 1551 20848
rect 0 20816 800 20846
rect 1485 20843 1551 20846
rect 4207 20704 4527 20705
rect 4207 20640 4215 20704
rect 4279 20640 4295 20704
rect 4359 20640 4375 20704
rect 4439 20640 4455 20704
rect 4519 20640 4527 20704
rect 4207 20639 4527 20640
rect 7471 20704 7791 20705
rect 7471 20640 7479 20704
rect 7543 20640 7559 20704
rect 7623 20640 7639 20704
rect 7703 20640 7719 20704
rect 7783 20640 7791 20704
rect 7471 20639 7791 20640
rect 9029 20634 9095 20637
rect 11200 20634 12000 20664
rect 9029 20632 12000 20634
rect 9029 20576 9034 20632
rect 9090 20576 12000 20632
rect 9029 20574 12000 20576
rect 9029 20571 9095 20574
rect 11200 20544 12000 20574
rect 0 20362 800 20392
rect 1485 20362 1551 20365
rect 0 20360 1551 20362
rect 0 20304 1490 20360
rect 1546 20304 1551 20360
rect 0 20302 1551 20304
rect 0 20272 800 20302
rect 1485 20299 1551 20302
rect 2576 20160 2896 20161
rect 2576 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2576 20095 2896 20096
rect 5839 20160 6159 20161
rect 5839 20096 5847 20160
rect 5911 20096 5927 20160
rect 5991 20096 6007 20160
rect 6071 20096 6087 20160
rect 6151 20096 6159 20160
rect 5839 20095 6159 20096
rect 9103 20160 9423 20161
rect 9103 20096 9111 20160
rect 9175 20096 9191 20160
rect 9255 20096 9271 20160
rect 9335 20096 9351 20160
rect 9415 20096 9423 20160
rect 9103 20095 9423 20096
rect 10133 19954 10199 19957
rect 11200 19954 12000 19984
rect 10133 19952 12000 19954
rect 10133 19896 10138 19952
rect 10194 19896 12000 19952
rect 10133 19894 12000 19896
rect 10133 19891 10199 19894
rect 11200 19864 12000 19894
rect 0 19682 800 19712
rect 1485 19682 1551 19685
rect 0 19680 1551 19682
rect 0 19624 1490 19680
rect 1546 19624 1551 19680
rect 0 19622 1551 19624
rect 0 19592 800 19622
rect 1485 19619 1551 19622
rect 4207 19616 4527 19617
rect 4207 19552 4215 19616
rect 4279 19552 4295 19616
rect 4359 19552 4375 19616
rect 4439 19552 4455 19616
rect 4519 19552 4527 19616
rect 4207 19551 4527 19552
rect 7471 19616 7791 19617
rect 7471 19552 7479 19616
rect 7543 19552 7559 19616
rect 7623 19552 7639 19616
rect 7703 19552 7719 19616
rect 7783 19552 7791 19616
rect 7471 19551 7791 19552
rect 0 19138 800 19168
rect 1485 19138 1551 19141
rect 0 19136 1551 19138
rect 0 19080 1490 19136
rect 1546 19080 1551 19136
rect 0 19078 1551 19080
rect 0 19048 800 19078
rect 1485 19075 1551 19078
rect 10225 19138 10291 19141
rect 11200 19138 12000 19168
rect 10225 19136 12000 19138
rect 10225 19080 10230 19136
rect 10286 19080 12000 19136
rect 10225 19078 12000 19080
rect 10225 19075 10291 19078
rect 2576 19072 2896 19073
rect 2576 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2576 19007 2896 19008
rect 5839 19072 6159 19073
rect 5839 19008 5847 19072
rect 5911 19008 5927 19072
rect 5991 19008 6007 19072
rect 6071 19008 6087 19072
rect 6151 19008 6159 19072
rect 5839 19007 6159 19008
rect 9103 19072 9423 19073
rect 9103 19008 9111 19072
rect 9175 19008 9191 19072
rect 9255 19008 9271 19072
rect 9335 19008 9351 19072
rect 9415 19008 9423 19072
rect 11200 19048 12000 19078
rect 9103 19007 9423 19008
rect 0 18594 800 18624
rect 1485 18594 1551 18597
rect 0 18592 1551 18594
rect 0 18536 1490 18592
rect 1546 18536 1551 18592
rect 0 18534 1551 18536
rect 0 18504 800 18534
rect 1485 18531 1551 18534
rect 4207 18528 4527 18529
rect 4207 18464 4215 18528
rect 4279 18464 4295 18528
rect 4359 18464 4375 18528
rect 4439 18464 4455 18528
rect 4519 18464 4527 18528
rect 4207 18463 4527 18464
rect 7471 18528 7791 18529
rect 7471 18464 7479 18528
rect 7543 18464 7559 18528
rect 7623 18464 7639 18528
rect 7703 18464 7719 18528
rect 7783 18464 7791 18528
rect 7471 18463 7791 18464
rect 11200 18368 12000 18488
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 2576 17984 2896 17985
rect 2576 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2576 17919 2896 17920
rect 5839 17984 6159 17985
rect 5839 17920 5847 17984
rect 5911 17920 5927 17984
rect 5991 17920 6007 17984
rect 6071 17920 6087 17984
rect 6151 17920 6159 17984
rect 5839 17919 6159 17920
rect 9103 17984 9423 17985
rect 9103 17920 9111 17984
rect 9175 17920 9191 17984
rect 9255 17920 9271 17984
rect 9335 17920 9351 17984
rect 9415 17920 9423 17984
rect 9103 17919 9423 17920
rect 11200 17552 12000 17672
rect 0 17506 800 17536
rect 1485 17506 1551 17509
rect 0 17504 1551 17506
rect 0 17448 1490 17504
rect 1546 17448 1551 17504
rect 0 17446 1551 17448
rect 0 17416 800 17446
rect 1485 17443 1551 17446
rect 4207 17440 4527 17441
rect 4207 17376 4215 17440
rect 4279 17376 4295 17440
rect 4359 17376 4375 17440
rect 4439 17376 4455 17440
rect 4519 17376 4527 17440
rect 4207 17375 4527 17376
rect 7471 17440 7791 17441
rect 7471 17376 7479 17440
rect 7543 17376 7559 17440
rect 7623 17376 7639 17440
rect 7703 17376 7719 17440
rect 7783 17376 7791 17440
rect 7471 17375 7791 17376
rect 0 16962 800 16992
rect 1485 16962 1551 16965
rect 0 16960 1551 16962
rect 0 16904 1490 16960
rect 1546 16904 1551 16960
rect 0 16902 1551 16904
rect 0 16872 800 16902
rect 1485 16899 1551 16902
rect 2576 16896 2896 16897
rect 2576 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2576 16831 2896 16832
rect 5839 16896 6159 16897
rect 5839 16832 5847 16896
rect 5911 16832 5927 16896
rect 5991 16832 6007 16896
rect 6071 16832 6087 16896
rect 6151 16832 6159 16896
rect 5839 16831 6159 16832
rect 9103 16896 9423 16897
rect 9103 16832 9111 16896
rect 9175 16832 9191 16896
rect 9255 16832 9271 16896
rect 9335 16832 9351 16896
rect 9415 16832 9423 16896
rect 11200 16872 12000 16992
rect 9103 16831 9423 16832
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 4207 16352 4527 16353
rect 4207 16288 4215 16352
rect 4279 16288 4295 16352
rect 4359 16288 4375 16352
rect 4439 16288 4455 16352
rect 4519 16288 4527 16352
rect 4207 16287 4527 16288
rect 7471 16352 7791 16353
rect 7471 16288 7479 16352
rect 7543 16288 7559 16352
rect 7623 16288 7639 16352
rect 7703 16288 7719 16352
rect 7783 16288 7791 16352
rect 7471 16287 7791 16288
rect 11200 16056 12000 16176
rect 0 15874 800 15904
rect 1485 15874 1551 15877
rect 0 15872 1551 15874
rect 0 15816 1490 15872
rect 1546 15816 1551 15872
rect 0 15814 1551 15816
rect 0 15784 800 15814
rect 1485 15811 1551 15814
rect 2576 15808 2896 15809
rect 2576 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2576 15743 2896 15744
rect 5839 15808 6159 15809
rect 5839 15744 5847 15808
rect 5911 15744 5927 15808
rect 5991 15744 6007 15808
rect 6071 15744 6087 15808
rect 6151 15744 6159 15808
rect 5839 15743 6159 15744
rect 9103 15808 9423 15809
rect 9103 15744 9111 15808
rect 9175 15744 9191 15808
rect 9255 15744 9271 15808
rect 9335 15744 9351 15808
rect 9415 15744 9423 15808
rect 9103 15743 9423 15744
rect 0 15330 800 15360
rect 1485 15330 1551 15333
rect 0 15328 1551 15330
rect 0 15272 1490 15328
rect 1546 15272 1551 15328
rect 0 15270 1551 15272
rect 0 15240 800 15270
rect 1485 15267 1551 15270
rect 4207 15264 4527 15265
rect 4207 15200 4215 15264
rect 4279 15200 4295 15264
rect 4359 15200 4375 15264
rect 4439 15200 4455 15264
rect 4519 15200 4527 15264
rect 4207 15199 4527 15200
rect 7471 15264 7791 15265
rect 7471 15200 7479 15264
rect 7543 15200 7559 15264
rect 7623 15200 7639 15264
rect 7703 15200 7719 15264
rect 7783 15200 7791 15264
rect 11200 15240 12000 15360
rect 7471 15199 7791 15200
rect 0 14786 800 14816
rect 1485 14786 1551 14789
rect 0 14784 1551 14786
rect 0 14728 1490 14784
rect 1546 14728 1551 14784
rect 0 14726 1551 14728
rect 0 14696 800 14726
rect 1485 14723 1551 14726
rect 2576 14720 2896 14721
rect 2576 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2576 14655 2896 14656
rect 5839 14720 6159 14721
rect 5839 14656 5847 14720
rect 5911 14656 5927 14720
rect 5991 14656 6007 14720
rect 6071 14656 6087 14720
rect 6151 14656 6159 14720
rect 5839 14655 6159 14656
rect 9103 14720 9423 14721
rect 9103 14656 9111 14720
rect 9175 14656 9191 14720
rect 9255 14656 9271 14720
rect 9335 14656 9351 14720
rect 9415 14656 9423 14720
rect 9103 14655 9423 14656
rect 11200 14560 12000 14680
rect 0 14242 800 14272
rect 1485 14242 1551 14245
rect 0 14240 1551 14242
rect 0 14184 1490 14240
rect 1546 14184 1551 14240
rect 0 14182 1551 14184
rect 0 14152 800 14182
rect 1485 14179 1551 14182
rect 4207 14176 4527 14177
rect 4207 14112 4215 14176
rect 4279 14112 4295 14176
rect 4359 14112 4375 14176
rect 4439 14112 4455 14176
rect 4519 14112 4527 14176
rect 4207 14111 4527 14112
rect 7471 14176 7791 14177
rect 7471 14112 7479 14176
rect 7543 14112 7559 14176
rect 7623 14112 7639 14176
rect 7703 14112 7719 14176
rect 7783 14112 7791 14176
rect 7471 14111 7791 14112
rect 11200 13744 12000 13864
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 2576 13632 2896 13633
rect 2576 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2576 13567 2896 13568
rect 5839 13632 6159 13633
rect 5839 13568 5847 13632
rect 5911 13568 5927 13632
rect 5991 13568 6007 13632
rect 6071 13568 6087 13632
rect 6151 13568 6159 13632
rect 5839 13567 6159 13568
rect 9103 13632 9423 13633
rect 9103 13568 9111 13632
rect 9175 13568 9191 13632
rect 9255 13568 9271 13632
rect 9335 13568 9351 13632
rect 9415 13568 9423 13632
rect 9103 13567 9423 13568
rect 4207 13088 4527 13089
rect 0 13018 800 13048
rect 4207 13024 4215 13088
rect 4279 13024 4295 13088
rect 4359 13024 4375 13088
rect 4439 13024 4455 13088
rect 4519 13024 4527 13088
rect 4207 13023 4527 13024
rect 7471 13088 7791 13089
rect 7471 13024 7479 13088
rect 7543 13024 7559 13088
rect 7623 13024 7639 13088
rect 7703 13024 7719 13088
rect 7783 13024 7791 13088
rect 11200 13064 12000 13184
rect 7471 13023 7791 13024
rect 1485 13018 1551 13021
rect 0 13016 1551 13018
rect 0 12960 1490 13016
rect 1546 12960 1551 13016
rect 0 12958 1551 12960
rect 0 12928 800 12958
rect 1485 12955 1551 12958
rect 2576 12544 2896 12545
rect 0 12474 800 12504
rect 2576 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2576 12479 2896 12480
rect 5839 12544 6159 12545
rect 5839 12480 5847 12544
rect 5911 12480 5927 12544
rect 5991 12480 6007 12544
rect 6071 12480 6087 12544
rect 6151 12480 6159 12544
rect 5839 12479 6159 12480
rect 9103 12544 9423 12545
rect 9103 12480 9111 12544
rect 9175 12480 9191 12544
rect 9255 12480 9271 12544
rect 9335 12480 9351 12544
rect 9415 12480 9423 12544
rect 9103 12479 9423 12480
rect 1485 12474 1551 12477
rect 0 12472 1551 12474
rect 0 12416 1490 12472
rect 1546 12416 1551 12472
rect 0 12414 1551 12416
rect 0 12384 800 12414
rect 1485 12411 1551 12414
rect 11200 12248 12000 12368
rect 4207 12000 4527 12001
rect 0 11930 800 11960
rect 4207 11936 4215 12000
rect 4279 11936 4295 12000
rect 4359 11936 4375 12000
rect 4439 11936 4455 12000
rect 4519 11936 4527 12000
rect 4207 11935 4527 11936
rect 7471 12000 7791 12001
rect 7471 11936 7479 12000
rect 7543 11936 7559 12000
rect 7623 11936 7639 12000
rect 7703 11936 7719 12000
rect 7783 11936 7791 12000
rect 7471 11935 7791 11936
rect 1485 11930 1551 11933
rect 0 11928 1551 11930
rect 0 11872 1490 11928
rect 1546 11872 1551 11928
rect 0 11870 1551 11872
rect 0 11840 800 11870
rect 1485 11867 1551 11870
rect 11200 11568 12000 11688
rect 2576 11456 2896 11457
rect 0 11386 800 11416
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 11391 2896 11392
rect 5839 11456 6159 11457
rect 5839 11392 5847 11456
rect 5911 11392 5927 11456
rect 5991 11392 6007 11456
rect 6071 11392 6087 11456
rect 6151 11392 6159 11456
rect 5839 11391 6159 11392
rect 9103 11456 9423 11457
rect 9103 11392 9111 11456
rect 9175 11392 9191 11456
rect 9255 11392 9271 11456
rect 9335 11392 9351 11456
rect 9415 11392 9423 11456
rect 9103 11391 9423 11392
rect 1485 11386 1551 11389
rect 0 11384 1551 11386
rect 0 11328 1490 11384
rect 1546 11328 1551 11384
rect 0 11326 1551 11328
rect 0 11296 800 11326
rect 1485 11323 1551 11326
rect 4207 10912 4527 10913
rect 0 10842 800 10872
rect 4207 10848 4215 10912
rect 4279 10848 4295 10912
rect 4359 10848 4375 10912
rect 4439 10848 4455 10912
rect 4519 10848 4527 10912
rect 4207 10847 4527 10848
rect 7471 10912 7791 10913
rect 7471 10848 7479 10912
rect 7543 10848 7559 10912
rect 7623 10848 7639 10912
rect 7703 10848 7719 10912
rect 7783 10848 7791 10912
rect 7471 10847 7791 10848
rect 1485 10842 1551 10845
rect 0 10840 1551 10842
rect 0 10784 1490 10840
rect 1546 10784 1551 10840
rect 0 10782 1551 10784
rect 0 10752 800 10782
rect 1485 10779 1551 10782
rect 11200 10752 12000 10872
rect 2576 10368 2896 10369
rect 0 10298 800 10328
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 10303 2896 10304
rect 5839 10368 6159 10369
rect 5839 10304 5847 10368
rect 5911 10304 5927 10368
rect 5991 10304 6007 10368
rect 6071 10304 6087 10368
rect 6151 10304 6159 10368
rect 5839 10303 6159 10304
rect 9103 10368 9423 10369
rect 9103 10304 9111 10368
rect 9175 10304 9191 10368
rect 9255 10304 9271 10368
rect 9335 10304 9351 10368
rect 9415 10304 9423 10368
rect 9103 10303 9423 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 11200 10072 12000 10192
rect 4207 9824 4527 9825
rect 0 9754 800 9784
rect 4207 9760 4215 9824
rect 4279 9760 4295 9824
rect 4359 9760 4375 9824
rect 4439 9760 4455 9824
rect 4519 9760 4527 9824
rect 4207 9759 4527 9760
rect 7471 9824 7791 9825
rect 7471 9760 7479 9824
rect 7543 9760 7559 9824
rect 7623 9760 7639 9824
rect 7703 9760 7719 9824
rect 7783 9760 7791 9824
rect 7471 9759 7791 9760
rect 1485 9754 1551 9757
rect 0 9752 1551 9754
rect 0 9696 1490 9752
rect 1546 9696 1551 9752
rect 0 9694 1551 9696
rect 0 9664 800 9694
rect 1485 9691 1551 9694
rect 2576 9280 2896 9281
rect 0 9210 800 9240
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 9215 2896 9216
rect 5839 9280 6159 9281
rect 5839 9216 5847 9280
rect 5911 9216 5927 9280
rect 5991 9216 6007 9280
rect 6071 9216 6087 9280
rect 6151 9216 6159 9280
rect 5839 9215 6159 9216
rect 9103 9280 9423 9281
rect 9103 9216 9111 9280
rect 9175 9216 9191 9280
rect 9255 9216 9271 9280
rect 9335 9216 9351 9280
rect 9415 9216 9423 9280
rect 11200 9256 12000 9376
rect 9103 9215 9423 9216
rect 2313 9210 2379 9213
rect 0 9208 2379 9210
rect 0 9152 2318 9208
rect 2374 9152 2379 9208
rect 0 9150 2379 9152
rect 0 9120 800 9150
rect 2313 9147 2379 9150
rect 4207 8736 4527 8737
rect 0 8666 800 8696
rect 4207 8672 4215 8736
rect 4279 8672 4295 8736
rect 4359 8672 4375 8736
rect 4439 8672 4455 8736
rect 4519 8672 4527 8736
rect 4207 8671 4527 8672
rect 7471 8736 7791 8737
rect 7471 8672 7479 8736
rect 7543 8672 7559 8736
rect 7623 8672 7639 8736
rect 7703 8672 7719 8736
rect 7783 8672 7791 8736
rect 7471 8671 7791 8672
rect 1485 8666 1551 8669
rect 0 8664 1551 8666
rect 0 8608 1490 8664
rect 1546 8608 1551 8664
rect 0 8606 1551 8608
rect 0 8576 800 8606
rect 1485 8603 1551 8606
rect 11200 8576 12000 8696
rect 2576 8192 2896 8193
rect 0 8122 800 8152
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 8127 2896 8128
rect 5839 8192 6159 8193
rect 5839 8128 5847 8192
rect 5911 8128 5927 8192
rect 5991 8128 6007 8192
rect 6071 8128 6087 8192
rect 6151 8128 6159 8192
rect 5839 8127 6159 8128
rect 9103 8192 9423 8193
rect 9103 8128 9111 8192
rect 9175 8128 9191 8192
rect 9255 8128 9271 8192
rect 9335 8128 9351 8192
rect 9415 8128 9423 8192
rect 9103 8127 9423 8128
rect 1393 8122 1459 8125
rect 0 8120 1459 8122
rect 0 8064 1398 8120
rect 1454 8064 1459 8120
rect 0 8062 1459 8064
rect 0 8032 800 8062
rect 1393 8059 1459 8062
rect 11200 7760 12000 7880
rect 4207 7648 4527 7649
rect 0 7578 800 7608
rect 4207 7584 4215 7648
rect 4279 7584 4295 7648
rect 4359 7584 4375 7648
rect 4439 7584 4455 7648
rect 4519 7584 4527 7648
rect 4207 7583 4527 7584
rect 7471 7648 7791 7649
rect 7471 7584 7479 7648
rect 7543 7584 7559 7648
rect 7623 7584 7639 7648
rect 7703 7584 7719 7648
rect 7783 7584 7791 7648
rect 7471 7583 7791 7584
rect 1485 7578 1551 7581
rect 0 7576 1551 7578
rect 0 7520 1490 7576
rect 1546 7520 1551 7576
rect 0 7518 1551 7520
rect 0 7488 800 7518
rect 1485 7515 1551 7518
rect 2576 7104 2896 7105
rect 0 7034 800 7064
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2576 7039 2896 7040
rect 5839 7104 6159 7105
rect 5839 7040 5847 7104
rect 5911 7040 5927 7104
rect 5991 7040 6007 7104
rect 6071 7040 6087 7104
rect 6151 7040 6159 7104
rect 5839 7039 6159 7040
rect 9103 7104 9423 7105
rect 9103 7040 9111 7104
rect 9175 7040 9191 7104
rect 9255 7040 9271 7104
rect 9335 7040 9351 7104
rect 9415 7040 9423 7104
rect 9103 7039 9423 7040
rect 2037 7034 2103 7037
rect 0 7032 2103 7034
rect 0 6976 2042 7032
rect 2098 6976 2103 7032
rect 0 6974 2103 6976
rect 0 6944 800 6974
rect 2037 6971 2103 6974
rect 11200 6944 12000 7064
rect 4207 6560 4527 6561
rect 4207 6496 4215 6560
rect 4279 6496 4295 6560
rect 4359 6496 4375 6560
rect 4439 6496 4455 6560
rect 4519 6496 4527 6560
rect 4207 6495 4527 6496
rect 7471 6560 7791 6561
rect 7471 6496 7479 6560
rect 7543 6496 7559 6560
rect 7623 6496 7639 6560
rect 7703 6496 7719 6560
rect 7783 6496 7791 6560
rect 7471 6495 7791 6496
rect 0 6354 800 6384
rect 1301 6354 1367 6357
rect 0 6352 1367 6354
rect 0 6296 1306 6352
rect 1362 6296 1367 6352
rect 0 6294 1367 6296
rect 0 6264 800 6294
rect 1301 6291 1367 6294
rect 10133 6354 10199 6357
rect 11200 6354 12000 6384
rect 10133 6352 12000 6354
rect 10133 6296 10138 6352
rect 10194 6296 12000 6352
rect 10133 6294 12000 6296
rect 10133 6291 10199 6294
rect 11200 6264 12000 6294
rect 2576 6016 2896 6017
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 5951 2896 5952
rect 5839 6016 6159 6017
rect 5839 5952 5847 6016
rect 5911 5952 5927 6016
rect 5991 5952 6007 6016
rect 6071 5952 6087 6016
rect 6151 5952 6159 6016
rect 5839 5951 6159 5952
rect 9103 6016 9423 6017
rect 9103 5952 9111 6016
rect 9175 5952 9191 6016
rect 9255 5952 9271 6016
rect 9335 5952 9351 6016
rect 9415 5952 9423 6016
rect 9103 5951 9423 5952
rect 0 5810 800 5840
rect 1485 5810 1551 5813
rect 0 5808 1551 5810
rect 0 5752 1490 5808
rect 1546 5752 1551 5808
rect 0 5750 1551 5752
rect 0 5720 800 5750
rect 1485 5747 1551 5750
rect 10133 5538 10199 5541
rect 11200 5538 12000 5568
rect 10133 5536 12000 5538
rect 10133 5480 10138 5536
rect 10194 5480 12000 5536
rect 10133 5478 12000 5480
rect 10133 5475 10199 5478
rect 4207 5472 4527 5473
rect 4207 5408 4215 5472
rect 4279 5408 4295 5472
rect 4359 5408 4375 5472
rect 4439 5408 4455 5472
rect 4519 5408 4527 5472
rect 4207 5407 4527 5408
rect 7471 5472 7791 5473
rect 7471 5408 7479 5472
rect 7543 5408 7559 5472
rect 7623 5408 7639 5472
rect 7703 5408 7719 5472
rect 7783 5408 7791 5472
rect 11200 5448 12000 5478
rect 7471 5407 7791 5408
rect 0 5266 800 5296
rect 1485 5266 1551 5269
rect 0 5264 1551 5266
rect 0 5208 1490 5264
rect 1546 5208 1551 5264
rect 0 5206 1551 5208
rect 0 5176 800 5206
rect 1485 5203 1551 5206
rect 2576 4928 2896 4929
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 4863 2896 4864
rect 5839 4928 6159 4929
rect 5839 4864 5847 4928
rect 5911 4864 5927 4928
rect 5991 4864 6007 4928
rect 6071 4864 6087 4928
rect 6151 4864 6159 4928
rect 5839 4863 6159 4864
rect 9103 4928 9423 4929
rect 9103 4864 9111 4928
rect 9175 4864 9191 4928
rect 9255 4864 9271 4928
rect 9335 4864 9351 4928
rect 9415 4864 9423 4928
rect 9103 4863 9423 4864
rect 10133 4858 10199 4861
rect 11200 4858 12000 4888
rect 10133 4856 12000 4858
rect 10133 4800 10138 4856
rect 10194 4800 12000 4856
rect 10133 4798 12000 4800
rect 10133 4795 10199 4798
rect 11200 4768 12000 4798
rect 0 4722 800 4752
rect 1485 4722 1551 4725
rect 0 4720 1551 4722
rect 0 4664 1490 4720
rect 1546 4664 1551 4720
rect 0 4662 1551 4664
rect 0 4632 800 4662
rect 1485 4659 1551 4662
rect 4207 4384 4527 4385
rect 4207 4320 4215 4384
rect 4279 4320 4295 4384
rect 4359 4320 4375 4384
rect 4439 4320 4455 4384
rect 4519 4320 4527 4384
rect 4207 4319 4527 4320
rect 7471 4384 7791 4385
rect 7471 4320 7479 4384
rect 7543 4320 7559 4384
rect 7623 4320 7639 4384
rect 7703 4320 7719 4384
rect 7783 4320 7791 4384
rect 7471 4319 7791 4320
rect 0 4178 800 4208
rect 1485 4178 1551 4181
rect 0 4176 1551 4178
rect 0 4120 1490 4176
rect 1546 4120 1551 4176
rect 0 4118 1551 4120
rect 0 4088 800 4118
rect 1485 4115 1551 4118
rect 10133 4042 10199 4045
rect 11200 4042 12000 4072
rect 10133 4040 12000 4042
rect 10133 3984 10138 4040
rect 10194 3984 12000 4040
rect 10133 3982 12000 3984
rect 10133 3979 10199 3982
rect 11200 3952 12000 3982
rect 2576 3840 2896 3841
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 3775 2896 3776
rect 5839 3840 6159 3841
rect 5839 3776 5847 3840
rect 5911 3776 5927 3840
rect 5991 3776 6007 3840
rect 6071 3776 6087 3840
rect 6151 3776 6159 3840
rect 5839 3775 6159 3776
rect 9103 3840 9423 3841
rect 9103 3776 9111 3840
rect 9175 3776 9191 3840
rect 9255 3776 9271 3840
rect 9335 3776 9351 3840
rect 9415 3776 9423 3840
rect 9103 3775 9423 3776
rect 0 3634 800 3664
rect 2313 3634 2379 3637
rect 0 3632 2379 3634
rect 0 3576 2318 3632
rect 2374 3576 2379 3632
rect 0 3574 2379 3576
rect 0 3544 800 3574
rect 2313 3571 2379 3574
rect 10133 3362 10199 3365
rect 11200 3362 12000 3392
rect 10133 3360 12000 3362
rect 10133 3304 10138 3360
rect 10194 3304 12000 3360
rect 10133 3302 12000 3304
rect 10133 3299 10199 3302
rect 4207 3296 4527 3297
rect 4207 3232 4215 3296
rect 4279 3232 4295 3296
rect 4359 3232 4375 3296
rect 4439 3232 4455 3296
rect 4519 3232 4527 3296
rect 4207 3231 4527 3232
rect 7471 3296 7791 3297
rect 7471 3232 7479 3296
rect 7543 3232 7559 3296
rect 7623 3232 7639 3296
rect 7703 3232 7719 3296
rect 7783 3232 7791 3296
rect 11200 3272 12000 3302
rect 7471 3231 7791 3232
rect 0 3090 800 3120
rect 1485 3090 1551 3093
rect 0 3088 1551 3090
rect 0 3032 1490 3088
rect 1546 3032 1551 3088
rect 0 3030 1551 3032
rect 0 3000 800 3030
rect 1485 3027 1551 3030
rect 2576 2752 2896 2753
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2687 2896 2688
rect 5839 2752 6159 2753
rect 5839 2688 5847 2752
rect 5911 2688 5927 2752
rect 5991 2688 6007 2752
rect 6071 2688 6087 2752
rect 6151 2688 6159 2752
rect 5839 2687 6159 2688
rect 9103 2752 9423 2753
rect 9103 2688 9111 2752
rect 9175 2688 9191 2752
rect 9255 2688 9271 2752
rect 9335 2688 9351 2752
rect 9415 2688 9423 2752
rect 9103 2687 9423 2688
rect 0 2546 800 2576
rect 1393 2546 1459 2549
rect 0 2544 1459 2546
rect 0 2488 1398 2544
rect 1454 2488 1459 2544
rect 0 2486 1459 2488
rect 0 2456 800 2486
rect 1393 2483 1459 2486
rect 10133 2546 10199 2549
rect 11200 2546 12000 2576
rect 10133 2544 12000 2546
rect 10133 2488 10138 2544
rect 10194 2488 12000 2544
rect 10133 2486 12000 2488
rect 10133 2483 10199 2486
rect 11200 2456 12000 2486
rect 4207 2208 4527 2209
rect 4207 2144 4215 2208
rect 4279 2144 4295 2208
rect 4359 2144 4375 2208
rect 4439 2144 4455 2208
rect 4519 2144 4527 2208
rect 4207 2143 4527 2144
rect 7471 2208 7791 2209
rect 7471 2144 7479 2208
rect 7543 2144 7559 2208
rect 7623 2144 7639 2208
rect 7703 2144 7719 2208
rect 7783 2144 7791 2208
rect 7471 2143 7791 2144
rect 0 2002 800 2032
rect 1485 2002 1551 2005
rect 0 2000 1551 2002
rect 0 1944 1490 2000
rect 1546 1944 1551 2000
rect 0 1942 1551 1944
rect 0 1912 800 1942
rect 1485 1939 1551 1942
rect 10133 1866 10199 1869
rect 11200 1866 12000 1896
rect 10133 1864 12000 1866
rect 10133 1808 10138 1864
rect 10194 1808 12000 1864
rect 10133 1806 12000 1808
rect 10133 1803 10199 1806
rect 11200 1776 12000 1806
rect 0 1458 800 1488
rect 3049 1458 3115 1461
rect 0 1456 3115 1458
rect 0 1400 3054 1456
rect 3110 1400 3115 1456
rect 0 1398 3115 1400
rect 0 1368 800 1398
rect 3049 1395 3115 1398
rect 11200 960 12000 1080
rect 0 914 800 944
rect 1393 914 1459 917
rect 0 912 1459 914
rect 0 856 1398 912
rect 1454 856 1459 912
rect 0 854 1459 856
rect 0 824 800 854
rect 1393 851 1459 854
rect 0 370 800 400
rect 2773 370 2839 373
rect 0 368 2839 370
rect 0 312 2778 368
rect 2834 312 2839 368
rect 0 310 2839 312
rect 0 280 800 310
rect 2773 307 2839 310
rect 11200 280 12000 400
<< via3 >>
rect 2584 77820 2648 77824
rect 2584 77764 2588 77820
rect 2588 77764 2644 77820
rect 2644 77764 2648 77820
rect 2584 77760 2648 77764
rect 2664 77820 2728 77824
rect 2664 77764 2668 77820
rect 2668 77764 2724 77820
rect 2724 77764 2728 77820
rect 2664 77760 2728 77764
rect 2744 77820 2808 77824
rect 2744 77764 2748 77820
rect 2748 77764 2804 77820
rect 2804 77764 2808 77820
rect 2744 77760 2808 77764
rect 2824 77820 2888 77824
rect 2824 77764 2828 77820
rect 2828 77764 2884 77820
rect 2884 77764 2888 77820
rect 2824 77760 2888 77764
rect 5847 77820 5911 77824
rect 5847 77764 5851 77820
rect 5851 77764 5907 77820
rect 5907 77764 5911 77820
rect 5847 77760 5911 77764
rect 5927 77820 5991 77824
rect 5927 77764 5931 77820
rect 5931 77764 5987 77820
rect 5987 77764 5991 77820
rect 5927 77760 5991 77764
rect 6007 77820 6071 77824
rect 6007 77764 6011 77820
rect 6011 77764 6067 77820
rect 6067 77764 6071 77820
rect 6007 77760 6071 77764
rect 6087 77820 6151 77824
rect 6087 77764 6091 77820
rect 6091 77764 6147 77820
rect 6147 77764 6151 77820
rect 6087 77760 6151 77764
rect 9111 77820 9175 77824
rect 9111 77764 9115 77820
rect 9115 77764 9171 77820
rect 9171 77764 9175 77820
rect 9111 77760 9175 77764
rect 9191 77820 9255 77824
rect 9191 77764 9195 77820
rect 9195 77764 9251 77820
rect 9251 77764 9255 77820
rect 9191 77760 9255 77764
rect 9271 77820 9335 77824
rect 9271 77764 9275 77820
rect 9275 77764 9331 77820
rect 9331 77764 9335 77820
rect 9271 77760 9335 77764
rect 9351 77820 9415 77824
rect 9351 77764 9355 77820
rect 9355 77764 9411 77820
rect 9411 77764 9415 77820
rect 9351 77760 9415 77764
rect 4215 77276 4279 77280
rect 4215 77220 4219 77276
rect 4219 77220 4275 77276
rect 4275 77220 4279 77276
rect 4215 77216 4279 77220
rect 4295 77276 4359 77280
rect 4295 77220 4299 77276
rect 4299 77220 4355 77276
rect 4355 77220 4359 77276
rect 4295 77216 4359 77220
rect 4375 77276 4439 77280
rect 4375 77220 4379 77276
rect 4379 77220 4435 77276
rect 4435 77220 4439 77276
rect 4375 77216 4439 77220
rect 4455 77276 4519 77280
rect 4455 77220 4459 77276
rect 4459 77220 4515 77276
rect 4515 77220 4519 77276
rect 4455 77216 4519 77220
rect 7479 77276 7543 77280
rect 7479 77220 7483 77276
rect 7483 77220 7539 77276
rect 7539 77220 7543 77276
rect 7479 77216 7543 77220
rect 7559 77276 7623 77280
rect 7559 77220 7563 77276
rect 7563 77220 7619 77276
rect 7619 77220 7623 77276
rect 7559 77216 7623 77220
rect 7639 77276 7703 77280
rect 7639 77220 7643 77276
rect 7643 77220 7699 77276
rect 7699 77220 7703 77276
rect 7639 77216 7703 77220
rect 7719 77276 7783 77280
rect 7719 77220 7723 77276
rect 7723 77220 7779 77276
rect 7779 77220 7783 77276
rect 7719 77216 7783 77220
rect 2584 76732 2648 76736
rect 2584 76676 2588 76732
rect 2588 76676 2644 76732
rect 2644 76676 2648 76732
rect 2584 76672 2648 76676
rect 2664 76732 2728 76736
rect 2664 76676 2668 76732
rect 2668 76676 2724 76732
rect 2724 76676 2728 76732
rect 2664 76672 2728 76676
rect 2744 76732 2808 76736
rect 2744 76676 2748 76732
rect 2748 76676 2804 76732
rect 2804 76676 2808 76732
rect 2744 76672 2808 76676
rect 2824 76732 2888 76736
rect 2824 76676 2828 76732
rect 2828 76676 2884 76732
rect 2884 76676 2888 76732
rect 2824 76672 2888 76676
rect 5847 76732 5911 76736
rect 5847 76676 5851 76732
rect 5851 76676 5907 76732
rect 5907 76676 5911 76732
rect 5847 76672 5911 76676
rect 5927 76732 5991 76736
rect 5927 76676 5931 76732
rect 5931 76676 5987 76732
rect 5987 76676 5991 76732
rect 5927 76672 5991 76676
rect 6007 76732 6071 76736
rect 6007 76676 6011 76732
rect 6011 76676 6067 76732
rect 6067 76676 6071 76732
rect 6007 76672 6071 76676
rect 6087 76732 6151 76736
rect 6087 76676 6091 76732
rect 6091 76676 6147 76732
rect 6147 76676 6151 76732
rect 6087 76672 6151 76676
rect 9111 76732 9175 76736
rect 9111 76676 9115 76732
rect 9115 76676 9171 76732
rect 9171 76676 9175 76732
rect 9111 76672 9175 76676
rect 9191 76732 9255 76736
rect 9191 76676 9195 76732
rect 9195 76676 9251 76732
rect 9251 76676 9255 76732
rect 9191 76672 9255 76676
rect 9271 76732 9335 76736
rect 9271 76676 9275 76732
rect 9275 76676 9331 76732
rect 9331 76676 9335 76732
rect 9271 76672 9335 76676
rect 9351 76732 9415 76736
rect 9351 76676 9355 76732
rect 9355 76676 9411 76732
rect 9411 76676 9415 76732
rect 9351 76672 9415 76676
rect 4215 76188 4279 76192
rect 4215 76132 4219 76188
rect 4219 76132 4275 76188
rect 4275 76132 4279 76188
rect 4215 76128 4279 76132
rect 4295 76188 4359 76192
rect 4295 76132 4299 76188
rect 4299 76132 4355 76188
rect 4355 76132 4359 76188
rect 4295 76128 4359 76132
rect 4375 76188 4439 76192
rect 4375 76132 4379 76188
rect 4379 76132 4435 76188
rect 4435 76132 4439 76188
rect 4375 76128 4439 76132
rect 4455 76188 4519 76192
rect 4455 76132 4459 76188
rect 4459 76132 4515 76188
rect 4515 76132 4519 76188
rect 4455 76128 4519 76132
rect 7479 76188 7543 76192
rect 7479 76132 7483 76188
rect 7483 76132 7539 76188
rect 7539 76132 7543 76188
rect 7479 76128 7543 76132
rect 7559 76188 7623 76192
rect 7559 76132 7563 76188
rect 7563 76132 7619 76188
rect 7619 76132 7623 76188
rect 7559 76128 7623 76132
rect 7639 76188 7703 76192
rect 7639 76132 7643 76188
rect 7643 76132 7699 76188
rect 7699 76132 7703 76188
rect 7639 76128 7703 76132
rect 7719 76188 7783 76192
rect 7719 76132 7723 76188
rect 7723 76132 7779 76188
rect 7779 76132 7783 76188
rect 7719 76128 7783 76132
rect 2584 75644 2648 75648
rect 2584 75588 2588 75644
rect 2588 75588 2644 75644
rect 2644 75588 2648 75644
rect 2584 75584 2648 75588
rect 2664 75644 2728 75648
rect 2664 75588 2668 75644
rect 2668 75588 2724 75644
rect 2724 75588 2728 75644
rect 2664 75584 2728 75588
rect 2744 75644 2808 75648
rect 2744 75588 2748 75644
rect 2748 75588 2804 75644
rect 2804 75588 2808 75644
rect 2744 75584 2808 75588
rect 2824 75644 2888 75648
rect 2824 75588 2828 75644
rect 2828 75588 2884 75644
rect 2884 75588 2888 75644
rect 2824 75584 2888 75588
rect 5847 75644 5911 75648
rect 5847 75588 5851 75644
rect 5851 75588 5907 75644
rect 5907 75588 5911 75644
rect 5847 75584 5911 75588
rect 5927 75644 5991 75648
rect 5927 75588 5931 75644
rect 5931 75588 5987 75644
rect 5987 75588 5991 75644
rect 5927 75584 5991 75588
rect 6007 75644 6071 75648
rect 6007 75588 6011 75644
rect 6011 75588 6067 75644
rect 6067 75588 6071 75644
rect 6007 75584 6071 75588
rect 6087 75644 6151 75648
rect 6087 75588 6091 75644
rect 6091 75588 6147 75644
rect 6147 75588 6151 75644
rect 6087 75584 6151 75588
rect 9111 75644 9175 75648
rect 9111 75588 9115 75644
rect 9115 75588 9171 75644
rect 9171 75588 9175 75644
rect 9111 75584 9175 75588
rect 9191 75644 9255 75648
rect 9191 75588 9195 75644
rect 9195 75588 9251 75644
rect 9251 75588 9255 75644
rect 9191 75584 9255 75588
rect 9271 75644 9335 75648
rect 9271 75588 9275 75644
rect 9275 75588 9331 75644
rect 9331 75588 9335 75644
rect 9271 75584 9335 75588
rect 9351 75644 9415 75648
rect 9351 75588 9355 75644
rect 9355 75588 9411 75644
rect 9411 75588 9415 75644
rect 9351 75584 9415 75588
rect 4215 75100 4279 75104
rect 4215 75044 4219 75100
rect 4219 75044 4275 75100
rect 4275 75044 4279 75100
rect 4215 75040 4279 75044
rect 4295 75100 4359 75104
rect 4295 75044 4299 75100
rect 4299 75044 4355 75100
rect 4355 75044 4359 75100
rect 4295 75040 4359 75044
rect 4375 75100 4439 75104
rect 4375 75044 4379 75100
rect 4379 75044 4435 75100
rect 4435 75044 4439 75100
rect 4375 75040 4439 75044
rect 4455 75100 4519 75104
rect 4455 75044 4459 75100
rect 4459 75044 4515 75100
rect 4515 75044 4519 75100
rect 4455 75040 4519 75044
rect 7479 75100 7543 75104
rect 7479 75044 7483 75100
rect 7483 75044 7539 75100
rect 7539 75044 7543 75100
rect 7479 75040 7543 75044
rect 7559 75100 7623 75104
rect 7559 75044 7563 75100
rect 7563 75044 7619 75100
rect 7619 75044 7623 75100
rect 7559 75040 7623 75044
rect 7639 75100 7703 75104
rect 7639 75044 7643 75100
rect 7643 75044 7699 75100
rect 7699 75044 7703 75100
rect 7639 75040 7703 75044
rect 7719 75100 7783 75104
rect 7719 75044 7723 75100
rect 7723 75044 7779 75100
rect 7779 75044 7783 75100
rect 7719 75040 7783 75044
rect 2584 74556 2648 74560
rect 2584 74500 2588 74556
rect 2588 74500 2644 74556
rect 2644 74500 2648 74556
rect 2584 74496 2648 74500
rect 2664 74556 2728 74560
rect 2664 74500 2668 74556
rect 2668 74500 2724 74556
rect 2724 74500 2728 74556
rect 2664 74496 2728 74500
rect 2744 74556 2808 74560
rect 2744 74500 2748 74556
rect 2748 74500 2804 74556
rect 2804 74500 2808 74556
rect 2744 74496 2808 74500
rect 2824 74556 2888 74560
rect 2824 74500 2828 74556
rect 2828 74500 2884 74556
rect 2884 74500 2888 74556
rect 2824 74496 2888 74500
rect 5847 74556 5911 74560
rect 5847 74500 5851 74556
rect 5851 74500 5907 74556
rect 5907 74500 5911 74556
rect 5847 74496 5911 74500
rect 5927 74556 5991 74560
rect 5927 74500 5931 74556
rect 5931 74500 5987 74556
rect 5987 74500 5991 74556
rect 5927 74496 5991 74500
rect 6007 74556 6071 74560
rect 6007 74500 6011 74556
rect 6011 74500 6067 74556
rect 6067 74500 6071 74556
rect 6007 74496 6071 74500
rect 6087 74556 6151 74560
rect 6087 74500 6091 74556
rect 6091 74500 6147 74556
rect 6147 74500 6151 74556
rect 6087 74496 6151 74500
rect 9111 74556 9175 74560
rect 9111 74500 9115 74556
rect 9115 74500 9171 74556
rect 9171 74500 9175 74556
rect 9111 74496 9175 74500
rect 9191 74556 9255 74560
rect 9191 74500 9195 74556
rect 9195 74500 9251 74556
rect 9251 74500 9255 74556
rect 9191 74496 9255 74500
rect 9271 74556 9335 74560
rect 9271 74500 9275 74556
rect 9275 74500 9331 74556
rect 9331 74500 9335 74556
rect 9271 74496 9335 74500
rect 9351 74556 9415 74560
rect 9351 74500 9355 74556
rect 9355 74500 9411 74556
rect 9411 74500 9415 74556
rect 9351 74496 9415 74500
rect 4215 74012 4279 74016
rect 4215 73956 4219 74012
rect 4219 73956 4275 74012
rect 4275 73956 4279 74012
rect 4215 73952 4279 73956
rect 4295 74012 4359 74016
rect 4295 73956 4299 74012
rect 4299 73956 4355 74012
rect 4355 73956 4359 74012
rect 4295 73952 4359 73956
rect 4375 74012 4439 74016
rect 4375 73956 4379 74012
rect 4379 73956 4435 74012
rect 4435 73956 4439 74012
rect 4375 73952 4439 73956
rect 4455 74012 4519 74016
rect 4455 73956 4459 74012
rect 4459 73956 4515 74012
rect 4515 73956 4519 74012
rect 4455 73952 4519 73956
rect 7479 74012 7543 74016
rect 7479 73956 7483 74012
rect 7483 73956 7539 74012
rect 7539 73956 7543 74012
rect 7479 73952 7543 73956
rect 7559 74012 7623 74016
rect 7559 73956 7563 74012
rect 7563 73956 7619 74012
rect 7619 73956 7623 74012
rect 7559 73952 7623 73956
rect 7639 74012 7703 74016
rect 7639 73956 7643 74012
rect 7643 73956 7699 74012
rect 7699 73956 7703 74012
rect 7639 73952 7703 73956
rect 7719 74012 7783 74016
rect 7719 73956 7723 74012
rect 7723 73956 7779 74012
rect 7779 73956 7783 74012
rect 7719 73952 7783 73956
rect 2584 73468 2648 73472
rect 2584 73412 2588 73468
rect 2588 73412 2644 73468
rect 2644 73412 2648 73468
rect 2584 73408 2648 73412
rect 2664 73468 2728 73472
rect 2664 73412 2668 73468
rect 2668 73412 2724 73468
rect 2724 73412 2728 73468
rect 2664 73408 2728 73412
rect 2744 73468 2808 73472
rect 2744 73412 2748 73468
rect 2748 73412 2804 73468
rect 2804 73412 2808 73468
rect 2744 73408 2808 73412
rect 2824 73468 2888 73472
rect 2824 73412 2828 73468
rect 2828 73412 2884 73468
rect 2884 73412 2888 73468
rect 2824 73408 2888 73412
rect 5847 73468 5911 73472
rect 5847 73412 5851 73468
rect 5851 73412 5907 73468
rect 5907 73412 5911 73468
rect 5847 73408 5911 73412
rect 5927 73468 5991 73472
rect 5927 73412 5931 73468
rect 5931 73412 5987 73468
rect 5987 73412 5991 73468
rect 5927 73408 5991 73412
rect 6007 73468 6071 73472
rect 6007 73412 6011 73468
rect 6011 73412 6067 73468
rect 6067 73412 6071 73468
rect 6007 73408 6071 73412
rect 6087 73468 6151 73472
rect 6087 73412 6091 73468
rect 6091 73412 6147 73468
rect 6147 73412 6151 73468
rect 6087 73408 6151 73412
rect 9111 73468 9175 73472
rect 9111 73412 9115 73468
rect 9115 73412 9171 73468
rect 9171 73412 9175 73468
rect 9111 73408 9175 73412
rect 9191 73468 9255 73472
rect 9191 73412 9195 73468
rect 9195 73412 9251 73468
rect 9251 73412 9255 73468
rect 9191 73408 9255 73412
rect 9271 73468 9335 73472
rect 9271 73412 9275 73468
rect 9275 73412 9331 73468
rect 9331 73412 9335 73468
rect 9271 73408 9335 73412
rect 9351 73468 9415 73472
rect 9351 73412 9355 73468
rect 9355 73412 9411 73468
rect 9411 73412 9415 73468
rect 9351 73408 9415 73412
rect 4215 72924 4279 72928
rect 4215 72868 4219 72924
rect 4219 72868 4275 72924
rect 4275 72868 4279 72924
rect 4215 72864 4279 72868
rect 4295 72924 4359 72928
rect 4295 72868 4299 72924
rect 4299 72868 4355 72924
rect 4355 72868 4359 72924
rect 4295 72864 4359 72868
rect 4375 72924 4439 72928
rect 4375 72868 4379 72924
rect 4379 72868 4435 72924
rect 4435 72868 4439 72924
rect 4375 72864 4439 72868
rect 4455 72924 4519 72928
rect 4455 72868 4459 72924
rect 4459 72868 4515 72924
rect 4515 72868 4519 72924
rect 4455 72864 4519 72868
rect 7479 72924 7543 72928
rect 7479 72868 7483 72924
rect 7483 72868 7539 72924
rect 7539 72868 7543 72924
rect 7479 72864 7543 72868
rect 7559 72924 7623 72928
rect 7559 72868 7563 72924
rect 7563 72868 7619 72924
rect 7619 72868 7623 72924
rect 7559 72864 7623 72868
rect 7639 72924 7703 72928
rect 7639 72868 7643 72924
rect 7643 72868 7699 72924
rect 7699 72868 7703 72924
rect 7639 72864 7703 72868
rect 7719 72924 7783 72928
rect 7719 72868 7723 72924
rect 7723 72868 7779 72924
rect 7779 72868 7783 72924
rect 7719 72864 7783 72868
rect 2584 72380 2648 72384
rect 2584 72324 2588 72380
rect 2588 72324 2644 72380
rect 2644 72324 2648 72380
rect 2584 72320 2648 72324
rect 2664 72380 2728 72384
rect 2664 72324 2668 72380
rect 2668 72324 2724 72380
rect 2724 72324 2728 72380
rect 2664 72320 2728 72324
rect 2744 72380 2808 72384
rect 2744 72324 2748 72380
rect 2748 72324 2804 72380
rect 2804 72324 2808 72380
rect 2744 72320 2808 72324
rect 2824 72380 2888 72384
rect 2824 72324 2828 72380
rect 2828 72324 2884 72380
rect 2884 72324 2888 72380
rect 2824 72320 2888 72324
rect 5847 72380 5911 72384
rect 5847 72324 5851 72380
rect 5851 72324 5907 72380
rect 5907 72324 5911 72380
rect 5847 72320 5911 72324
rect 5927 72380 5991 72384
rect 5927 72324 5931 72380
rect 5931 72324 5987 72380
rect 5987 72324 5991 72380
rect 5927 72320 5991 72324
rect 6007 72380 6071 72384
rect 6007 72324 6011 72380
rect 6011 72324 6067 72380
rect 6067 72324 6071 72380
rect 6007 72320 6071 72324
rect 6087 72380 6151 72384
rect 6087 72324 6091 72380
rect 6091 72324 6147 72380
rect 6147 72324 6151 72380
rect 6087 72320 6151 72324
rect 9111 72380 9175 72384
rect 9111 72324 9115 72380
rect 9115 72324 9171 72380
rect 9171 72324 9175 72380
rect 9111 72320 9175 72324
rect 9191 72380 9255 72384
rect 9191 72324 9195 72380
rect 9195 72324 9251 72380
rect 9251 72324 9255 72380
rect 9191 72320 9255 72324
rect 9271 72380 9335 72384
rect 9271 72324 9275 72380
rect 9275 72324 9331 72380
rect 9331 72324 9335 72380
rect 9271 72320 9335 72324
rect 9351 72380 9415 72384
rect 9351 72324 9355 72380
rect 9355 72324 9411 72380
rect 9411 72324 9415 72380
rect 9351 72320 9415 72324
rect 4215 71836 4279 71840
rect 4215 71780 4219 71836
rect 4219 71780 4275 71836
rect 4275 71780 4279 71836
rect 4215 71776 4279 71780
rect 4295 71836 4359 71840
rect 4295 71780 4299 71836
rect 4299 71780 4355 71836
rect 4355 71780 4359 71836
rect 4295 71776 4359 71780
rect 4375 71836 4439 71840
rect 4375 71780 4379 71836
rect 4379 71780 4435 71836
rect 4435 71780 4439 71836
rect 4375 71776 4439 71780
rect 4455 71836 4519 71840
rect 4455 71780 4459 71836
rect 4459 71780 4515 71836
rect 4515 71780 4519 71836
rect 4455 71776 4519 71780
rect 7479 71836 7543 71840
rect 7479 71780 7483 71836
rect 7483 71780 7539 71836
rect 7539 71780 7543 71836
rect 7479 71776 7543 71780
rect 7559 71836 7623 71840
rect 7559 71780 7563 71836
rect 7563 71780 7619 71836
rect 7619 71780 7623 71836
rect 7559 71776 7623 71780
rect 7639 71836 7703 71840
rect 7639 71780 7643 71836
rect 7643 71780 7699 71836
rect 7699 71780 7703 71836
rect 7639 71776 7703 71780
rect 7719 71836 7783 71840
rect 7719 71780 7723 71836
rect 7723 71780 7779 71836
rect 7779 71780 7783 71836
rect 7719 71776 7783 71780
rect 2584 71292 2648 71296
rect 2584 71236 2588 71292
rect 2588 71236 2644 71292
rect 2644 71236 2648 71292
rect 2584 71232 2648 71236
rect 2664 71292 2728 71296
rect 2664 71236 2668 71292
rect 2668 71236 2724 71292
rect 2724 71236 2728 71292
rect 2664 71232 2728 71236
rect 2744 71292 2808 71296
rect 2744 71236 2748 71292
rect 2748 71236 2804 71292
rect 2804 71236 2808 71292
rect 2744 71232 2808 71236
rect 2824 71292 2888 71296
rect 2824 71236 2828 71292
rect 2828 71236 2884 71292
rect 2884 71236 2888 71292
rect 2824 71232 2888 71236
rect 5847 71292 5911 71296
rect 5847 71236 5851 71292
rect 5851 71236 5907 71292
rect 5907 71236 5911 71292
rect 5847 71232 5911 71236
rect 5927 71292 5991 71296
rect 5927 71236 5931 71292
rect 5931 71236 5987 71292
rect 5987 71236 5991 71292
rect 5927 71232 5991 71236
rect 6007 71292 6071 71296
rect 6007 71236 6011 71292
rect 6011 71236 6067 71292
rect 6067 71236 6071 71292
rect 6007 71232 6071 71236
rect 6087 71292 6151 71296
rect 6087 71236 6091 71292
rect 6091 71236 6147 71292
rect 6147 71236 6151 71292
rect 6087 71232 6151 71236
rect 9111 71292 9175 71296
rect 9111 71236 9115 71292
rect 9115 71236 9171 71292
rect 9171 71236 9175 71292
rect 9111 71232 9175 71236
rect 9191 71292 9255 71296
rect 9191 71236 9195 71292
rect 9195 71236 9251 71292
rect 9251 71236 9255 71292
rect 9191 71232 9255 71236
rect 9271 71292 9335 71296
rect 9271 71236 9275 71292
rect 9275 71236 9331 71292
rect 9331 71236 9335 71292
rect 9271 71232 9335 71236
rect 9351 71292 9415 71296
rect 9351 71236 9355 71292
rect 9355 71236 9411 71292
rect 9411 71236 9415 71292
rect 9351 71232 9415 71236
rect 4215 70748 4279 70752
rect 4215 70692 4219 70748
rect 4219 70692 4275 70748
rect 4275 70692 4279 70748
rect 4215 70688 4279 70692
rect 4295 70748 4359 70752
rect 4295 70692 4299 70748
rect 4299 70692 4355 70748
rect 4355 70692 4359 70748
rect 4295 70688 4359 70692
rect 4375 70748 4439 70752
rect 4375 70692 4379 70748
rect 4379 70692 4435 70748
rect 4435 70692 4439 70748
rect 4375 70688 4439 70692
rect 4455 70748 4519 70752
rect 4455 70692 4459 70748
rect 4459 70692 4515 70748
rect 4515 70692 4519 70748
rect 4455 70688 4519 70692
rect 7479 70748 7543 70752
rect 7479 70692 7483 70748
rect 7483 70692 7539 70748
rect 7539 70692 7543 70748
rect 7479 70688 7543 70692
rect 7559 70748 7623 70752
rect 7559 70692 7563 70748
rect 7563 70692 7619 70748
rect 7619 70692 7623 70748
rect 7559 70688 7623 70692
rect 7639 70748 7703 70752
rect 7639 70692 7643 70748
rect 7643 70692 7699 70748
rect 7699 70692 7703 70748
rect 7639 70688 7703 70692
rect 7719 70748 7783 70752
rect 7719 70692 7723 70748
rect 7723 70692 7779 70748
rect 7779 70692 7783 70748
rect 7719 70688 7783 70692
rect 2584 70204 2648 70208
rect 2584 70148 2588 70204
rect 2588 70148 2644 70204
rect 2644 70148 2648 70204
rect 2584 70144 2648 70148
rect 2664 70204 2728 70208
rect 2664 70148 2668 70204
rect 2668 70148 2724 70204
rect 2724 70148 2728 70204
rect 2664 70144 2728 70148
rect 2744 70204 2808 70208
rect 2744 70148 2748 70204
rect 2748 70148 2804 70204
rect 2804 70148 2808 70204
rect 2744 70144 2808 70148
rect 2824 70204 2888 70208
rect 2824 70148 2828 70204
rect 2828 70148 2884 70204
rect 2884 70148 2888 70204
rect 2824 70144 2888 70148
rect 5847 70204 5911 70208
rect 5847 70148 5851 70204
rect 5851 70148 5907 70204
rect 5907 70148 5911 70204
rect 5847 70144 5911 70148
rect 5927 70204 5991 70208
rect 5927 70148 5931 70204
rect 5931 70148 5987 70204
rect 5987 70148 5991 70204
rect 5927 70144 5991 70148
rect 6007 70204 6071 70208
rect 6007 70148 6011 70204
rect 6011 70148 6067 70204
rect 6067 70148 6071 70204
rect 6007 70144 6071 70148
rect 6087 70204 6151 70208
rect 6087 70148 6091 70204
rect 6091 70148 6147 70204
rect 6147 70148 6151 70204
rect 6087 70144 6151 70148
rect 9111 70204 9175 70208
rect 9111 70148 9115 70204
rect 9115 70148 9171 70204
rect 9171 70148 9175 70204
rect 9111 70144 9175 70148
rect 9191 70204 9255 70208
rect 9191 70148 9195 70204
rect 9195 70148 9251 70204
rect 9251 70148 9255 70204
rect 9191 70144 9255 70148
rect 9271 70204 9335 70208
rect 9271 70148 9275 70204
rect 9275 70148 9331 70204
rect 9331 70148 9335 70204
rect 9271 70144 9335 70148
rect 9351 70204 9415 70208
rect 9351 70148 9355 70204
rect 9355 70148 9411 70204
rect 9411 70148 9415 70204
rect 9351 70144 9415 70148
rect 4215 69660 4279 69664
rect 4215 69604 4219 69660
rect 4219 69604 4275 69660
rect 4275 69604 4279 69660
rect 4215 69600 4279 69604
rect 4295 69660 4359 69664
rect 4295 69604 4299 69660
rect 4299 69604 4355 69660
rect 4355 69604 4359 69660
rect 4295 69600 4359 69604
rect 4375 69660 4439 69664
rect 4375 69604 4379 69660
rect 4379 69604 4435 69660
rect 4435 69604 4439 69660
rect 4375 69600 4439 69604
rect 4455 69660 4519 69664
rect 4455 69604 4459 69660
rect 4459 69604 4515 69660
rect 4515 69604 4519 69660
rect 4455 69600 4519 69604
rect 7479 69660 7543 69664
rect 7479 69604 7483 69660
rect 7483 69604 7539 69660
rect 7539 69604 7543 69660
rect 7479 69600 7543 69604
rect 7559 69660 7623 69664
rect 7559 69604 7563 69660
rect 7563 69604 7619 69660
rect 7619 69604 7623 69660
rect 7559 69600 7623 69604
rect 7639 69660 7703 69664
rect 7639 69604 7643 69660
rect 7643 69604 7699 69660
rect 7699 69604 7703 69660
rect 7639 69600 7703 69604
rect 7719 69660 7783 69664
rect 7719 69604 7723 69660
rect 7723 69604 7779 69660
rect 7779 69604 7783 69660
rect 7719 69600 7783 69604
rect 2584 69116 2648 69120
rect 2584 69060 2588 69116
rect 2588 69060 2644 69116
rect 2644 69060 2648 69116
rect 2584 69056 2648 69060
rect 2664 69116 2728 69120
rect 2664 69060 2668 69116
rect 2668 69060 2724 69116
rect 2724 69060 2728 69116
rect 2664 69056 2728 69060
rect 2744 69116 2808 69120
rect 2744 69060 2748 69116
rect 2748 69060 2804 69116
rect 2804 69060 2808 69116
rect 2744 69056 2808 69060
rect 2824 69116 2888 69120
rect 2824 69060 2828 69116
rect 2828 69060 2884 69116
rect 2884 69060 2888 69116
rect 2824 69056 2888 69060
rect 5847 69116 5911 69120
rect 5847 69060 5851 69116
rect 5851 69060 5907 69116
rect 5907 69060 5911 69116
rect 5847 69056 5911 69060
rect 5927 69116 5991 69120
rect 5927 69060 5931 69116
rect 5931 69060 5987 69116
rect 5987 69060 5991 69116
rect 5927 69056 5991 69060
rect 6007 69116 6071 69120
rect 6007 69060 6011 69116
rect 6011 69060 6067 69116
rect 6067 69060 6071 69116
rect 6007 69056 6071 69060
rect 6087 69116 6151 69120
rect 6087 69060 6091 69116
rect 6091 69060 6147 69116
rect 6147 69060 6151 69116
rect 6087 69056 6151 69060
rect 9111 69116 9175 69120
rect 9111 69060 9115 69116
rect 9115 69060 9171 69116
rect 9171 69060 9175 69116
rect 9111 69056 9175 69060
rect 9191 69116 9255 69120
rect 9191 69060 9195 69116
rect 9195 69060 9251 69116
rect 9251 69060 9255 69116
rect 9191 69056 9255 69060
rect 9271 69116 9335 69120
rect 9271 69060 9275 69116
rect 9275 69060 9331 69116
rect 9331 69060 9335 69116
rect 9271 69056 9335 69060
rect 9351 69116 9415 69120
rect 9351 69060 9355 69116
rect 9355 69060 9411 69116
rect 9411 69060 9415 69116
rect 9351 69056 9415 69060
rect 4215 68572 4279 68576
rect 4215 68516 4219 68572
rect 4219 68516 4275 68572
rect 4275 68516 4279 68572
rect 4215 68512 4279 68516
rect 4295 68572 4359 68576
rect 4295 68516 4299 68572
rect 4299 68516 4355 68572
rect 4355 68516 4359 68572
rect 4295 68512 4359 68516
rect 4375 68572 4439 68576
rect 4375 68516 4379 68572
rect 4379 68516 4435 68572
rect 4435 68516 4439 68572
rect 4375 68512 4439 68516
rect 4455 68572 4519 68576
rect 4455 68516 4459 68572
rect 4459 68516 4515 68572
rect 4515 68516 4519 68572
rect 4455 68512 4519 68516
rect 7479 68572 7543 68576
rect 7479 68516 7483 68572
rect 7483 68516 7539 68572
rect 7539 68516 7543 68572
rect 7479 68512 7543 68516
rect 7559 68572 7623 68576
rect 7559 68516 7563 68572
rect 7563 68516 7619 68572
rect 7619 68516 7623 68572
rect 7559 68512 7623 68516
rect 7639 68572 7703 68576
rect 7639 68516 7643 68572
rect 7643 68516 7699 68572
rect 7699 68516 7703 68572
rect 7639 68512 7703 68516
rect 7719 68572 7783 68576
rect 7719 68516 7723 68572
rect 7723 68516 7779 68572
rect 7779 68516 7783 68572
rect 7719 68512 7783 68516
rect 2584 68028 2648 68032
rect 2584 67972 2588 68028
rect 2588 67972 2644 68028
rect 2644 67972 2648 68028
rect 2584 67968 2648 67972
rect 2664 68028 2728 68032
rect 2664 67972 2668 68028
rect 2668 67972 2724 68028
rect 2724 67972 2728 68028
rect 2664 67968 2728 67972
rect 2744 68028 2808 68032
rect 2744 67972 2748 68028
rect 2748 67972 2804 68028
rect 2804 67972 2808 68028
rect 2744 67968 2808 67972
rect 2824 68028 2888 68032
rect 2824 67972 2828 68028
rect 2828 67972 2884 68028
rect 2884 67972 2888 68028
rect 2824 67968 2888 67972
rect 5847 68028 5911 68032
rect 5847 67972 5851 68028
rect 5851 67972 5907 68028
rect 5907 67972 5911 68028
rect 5847 67968 5911 67972
rect 5927 68028 5991 68032
rect 5927 67972 5931 68028
rect 5931 67972 5987 68028
rect 5987 67972 5991 68028
rect 5927 67968 5991 67972
rect 6007 68028 6071 68032
rect 6007 67972 6011 68028
rect 6011 67972 6067 68028
rect 6067 67972 6071 68028
rect 6007 67968 6071 67972
rect 6087 68028 6151 68032
rect 6087 67972 6091 68028
rect 6091 67972 6147 68028
rect 6147 67972 6151 68028
rect 6087 67968 6151 67972
rect 9111 68028 9175 68032
rect 9111 67972 9115 68028
rect 9115 67972 9171 68028
rect 9171 67972 9175 68028
rect 9111 67968 9175 67972
rect 9191 68028 9255 68032
rect 9191 67972 9195 68028
rect 9195 67972 9251 68028
rect 9251 67972 9255 68028
rect 9191 67968 9255 67972
rect 9271 68028 9335 68032
rect 9271 67972 9275 68028
rect 9275 67972 9331 68028
rect 9331 67972 9335 68028
rect 9271 67968 9335 67972
rect 9351 68028 9415 68032
rect 9351 67972 9355 68028
rect 9355 67972 9411 68028
rect 9411 67972 9415 68028
rect 9351 67968 9415 67972
rect 4215 67484 4279 67488
rect 4215 67428 4219 67484
rect 4219 67428 4275 67484
rect 4275 67428 4279 67484
rect 4215 67424 4279 67428
rect 4295 67484 4359 67488
rect 4295 67428 4299 67484
rect 4299 67428 4355 67484
rect 4355 67428 4359 67484
rect 4295 67424 4359 67428
rect 4375 67484 4439 67488
rect 4375 67428 4379 67484
rect 4379 67428 4435 67484
rect 4435 67428 4439 67484
rect 4375 67424 4439 67428
rect 4455 67484 4519 67488
rect 4455 67428 4459 67484
rect 4459 67428 4515 67484
rect 4515 67428 4519 67484
rect 4455 67424 4519 67428
rect 7479 67484 7543 67488
rect 7479 67428 7483 67484
rect 7483 67428 7539 67484
rect 7539 67428 7543 67484
rect 7479 67424 7543 67428
rect 7559 67484 7623 67488
rect 7559 67428 7563 67484
rect 7563 67428 7619 67484
rect 7619 67428 7623 67484
rect 7559 67424 7623 67428
rect 7639 67484 7703 67488
rect 7639 67428 7643 67484
rect 7643 67428 7699 67484
rect 7699 67428 7703 67484
rect 7639 67424 7703 67428
rect 7719 67484 7783 67488
rect 7719 67428 7723 67484
rect 7723 67428 7779 67484
rect 7779 67428 7783 67484
rect 7719 67424 7783 67428
rect 2584 66940 2648 66944
rect 2584 66884 2588 66940
rect 2588 66884 2644 66940
rect 2644 66884 2648 66940
rect 2584 66880 2648 66884
rect 2664 66940 2728 66944
rect 2664 66884 2668 66940
rect 2668 66884 2724 66940
rect 2724 66884 2728 66940
rect 2664 66880 2728 66884
rect 2744 66940 2808 66944
rect 2744 66884 2748 66940
rect 2748 66884 2804 66940
rect 2804 66884 2808 66940
rect 2744 66880 2808 66884
rect 2824 66940 2888 66944
rect 2824 66884 2828 66940
rect 2828 66884 2884 66940
rect 2884 66884 2888 66940
rect 2824 66880 2888 66884
rect 5847 66940 5911 66944
rect 5847 66884 5851 66940
rect 5851 66884 5907 66940
rect 5907 66884 5911 66940
rect 5847 66880 5911 66884
rect 5927 66940 5991 66944
rect 5927 66884 5931 66940
rect 5931 66884 5987 66940
rect 5987 66884 5991 66940
rect 5927 66880 5991 66884
rect 6007 66940 6071 66944
rect 6007 66884 6011 66940
rect 6011 66884 6067 66940
rect 6067 66884 6071 66940
rect 6007 66880 6071 66884
rect 6087 66940 6151 66944
rect 6087 66884 6091 66940
rect 6091 66884 6147 66940
rect 6147 66884 6151 66940
rect 6087 66880 6151 66884
rect 9111 66940 9175 66944
rect 9111 66884 9115 66940
rect 9115 66884 9171 66940
rect 9171 66884 9175 66940
rect 9111 66880 9175 66884
rect 9191 66940 9255 66944
rect 9191 66884 9195 66940
rect 9195 66884 9251 66940
rect 9251 66884 9255 66940
rect 9191 66880 9255 66884
rect 9271 66940 9335 66944
rect 9271 66884 9275 66940
rect 9275 66884 9331 66940
rect 9331 66884 9335 66940
rect 9271 66880 9335 66884
rect 9351 66940 9415 66944
rect 9351 66884 9355 66940
rect 9355 66884 9411 66940
rect 9411 66884 9415 66940
rect 9351 66880 9415 66884
rect 4215 66396 4279 66400
rect 4215 66340 4219 66396
rect 4219 66340 4275 66396
rect 4275 66340 4279 66396
rect 4215 66336 4279 66340
rect 4295 66396 4359 66400
rect 4295 66340 4299 66396
rect 4299 66340 4355 66396
rect 4355 66340 4359 66396
rect 4295 66336 4359 66340
rect 4375 66396 4439 66400
rect 4375 66340 4379 66396
rect 4379 66340 4435 66396
rect 4435 66340 4439 66396
rect 4375 66336 4439 66340
rect 4455 66396 4519 66400
rect 4455 66340 4459 66396
rect 4459 66340 4515 66396
rect 4515 66340 4519 66396
rect 4455 66336 4519 66340
rect 7479 66396 7543 66400
rect 7479 66340 7483 66396
rect 7483 66340 7539 66396
rect 7539 66340 7543 66396
rect 7479 66336 7543 66340
rect 7559 66396 7623 66400
rect 7559 66340 7563 66396
rect 7563 66340 7619 66396
rect 7619 66340 7623 66396
rect 7559 66336 7623 66340
rect 7639 66396 7703 66400
rect 7639 66340 7643 66396
rect 7643 66340 7699 66396
rect 7699 66340 7703 66396
rect 7639 66336 7703 66340
rect 7719 66396 7783 66400
rect 7719 66340 7723 66396
rect 7723 66340 7779 66396
rect 7779 66340 7783 66396
rect 7719 66336 7783 66340
rect 2584 65852 2648 65856
rect 2584 65796 2588 65852
rect 2588 65796 2644 65852
rect 2644 65796 2648 65852
rect 2584 65792 2648 65796
rect 2664 65852 2728 65856
rect 2664 65796 2668 65852
rect 2668 65796 2724 65852
rect 2724 65796 2728 65852
rect 2664 65792 2728 65796
rect 2744 65852 2808 65856
rect 2744 65796 2748 65852
rect 2748 65796 2804 65852
rect 2804 65796 2808 65852
rect 2744 65792 2808 65796
rect 2824 65852 2888 65856
rect 2824 65796 2828 65852
rect 2828 65796 2884 65852
rect 2884 65796 2888 65852
rect 2824 65792 2888 65796
rect 5847 65852 5911 65856
rect 5847 65796 5851 65852
rect 5851 65796 5907 65852
rect 5907 65796 5911 65852
rect 5847 65792 5911 65796
rect 5927 65852 5991 65856
rect 5927 65796 5931 65852
rect 5931 65796 5987 65852
rect 5987 65796 5991 65852
rect 5927 65792 5991 65796
rect 6007 65852 6071 65856
rect 6007 65796 6011 65852
rect 6011 65796 6067 65852
rect 6067 65796 6071 65852
rect 6007 65792 6071 65796
rect 6087 65852 6151 65856
rect 6087 65796 6091 65852
rect 6091 65796 6147 65852
rect 6147 65796 6151 65852
rect 6087 65792 6151 65796
rect 9111 65852 9175 65856
rect 9111 65796 9115 65852
rect 9115 65796 9171 65852
rect 9171 65796 9175 65852
rect 9111 65792 9175 65796
rect 9191 65852 9255 65856
rect 9191 65796 9195 65852
rect 9195 65796 9251 65852
rect 9251 65796 9255 65852
rect 9191 65792 9255 65796
rect 9271 65852 9335 65856
rect 9271 65796 9275 65852
rect 9275 65796 9331 65852
rect 9331 65796 9335 65852
rect 9271 65792 9335 65796
rect 9351 65852 9415 65856
rect 9351 65796 9355 65852
rect 9355 65796 9411 65852
rect 9411 65796 9415 65852
rect 9351 65792 9415 65796
rect 4215 65308 4279 65312
rect 4215 65252 4219 65308
rect 4219 65252 4275 65308
rect 4275 65252 4279 65308
rect 4215 65248 4279 65252
rect 4295 65308 4359 65312
rect 4295 65252 4299 65308
rect 4299 65252 4355 65308
rect 4355 65252 4359 65308
rect 4295 65248 4359 65252
rect 4375 65308 4439 65312
rect 4375 65252 4379 65308
rect 4379 65252 4435 65308
rect 4435 65252 4439 65308
rect 4375 65248 4439 65252
rect 4455 65308 4519 65312
rect 4455 65252 4459 65308
rect 4459 65252 4515 65308
rect 4515 65252 4519 65308
rect 4455 65248 4519 65252
rect 7479 65308 7543 65312
rect 7479 65252 7483 65308
rect 7483 65252 7539 65308
rect 7539 65252 7543 65308
rect 7479 65248 7543 65252
rect 7559 65308 7623 65312
rect 7559 65252 7563 65308
rect 7563 65252 7619 65308
rect 7619 65252 7623 65308
rect 7559 65248 7623 65252
rect 7639 65308 7703 65312
rect 7639 65252 7643 65308
rect 7643 65252 7699 65308
rect 7699 65252 7703 65308
rect 7639 65248 7703 65252
rect 7719 65308 7783 65312
rect 7719 65252 7723 65308
rect 7723 65252 7779 65308
rect 7779 65252 7783 65308
rect 7719 65248 7783 65252
rect 2584 64764 2648 64768
rect 2584 64708 2588 64764
rect 2588 64708 2644 64764
rect 2644 64708 2648 64764
rect 2584 64704 2648 64708
rect 2664 64764 2728 64768
rect 2664 64708 2668 64764
rect 2668 64708 2724 64764
rect 2724 64708 2728 64764
rect 2664 64704 2728 64708
rect 2744 64764 2808 64768
rect 2744 64708 2748 64764
rect 2748 64708 2804 64764
rect 2804 64708 2808 64764
rect 2744 64704 2808 64708
rect 2824 64764 2888 64768
rect 2824 64708 2828 64764
rect 2828 64708 2884 64764
rect 2884 64708 2888 64764
rect 2824 64704 2888 64708
rect 5847 64764 5911 64768
rect 5847 64708 5851 64764
rect 5851 64708 5907 64764
rect 5907 64708 5911 64764
rect 5847 64704 5911 64708
rect 5927 64764 5991 64768
rect 5927 64708 5931 64764
rect 5931 64708 5987 64764
rect 5987 64708 5991 64764
rect 5927 64704 5991 64708
rect 6007 64764 6071 64768
rect 6007 64708 6011 64764
rect 6011 64708 6067 64764
rect 6067 64708 6071 64764
rect 6007 64704 6071 64708
rect 6087 64764 6151 64768
rect 6087 64708 6091 64764
rect 6091 64708 6147 64764
rect 6147 64708 6151 64764
rect 6087 64704 6151 64708
rect 9111 64764 9175 64768
rect 9111 64708 9115 64764
rect 9115 64708 9171 64764
rect 9171 64708 9175 64764
rect 9111 64704 9175 64708
rect 9191 64764 9255 64768
rect 9191 64708 9195 64764
rect 9195 64708 9251 64764
rect 9251 64708 9255 64764
rect 9191 64704 9255 64708
rect 9271 64764 9335 64768
rect 9271 64708 9275 64764
rect 9275 64708 9331 64764
rect 9331 64708 9335 64764
rect 9271 64704 9335 64708
rect 9351 64764 9415 64768
rect 9351 64708 9355 64764
rect 9355 64708 9411 64764
rect 9411 64708 9415 64764
rect 9351 64704 9415 64708
rect 4215 64220 4279 64224
rect 4215 64164 4219 64220
rect 4219 64164 4275 64220
rect 4275 64164 4279 64220
rect 4215 64160 4279 64164
rect 4295 64220 4359 64224
rect 4295 64164 4299 64220
rect 4299 64164 4355 64220
rect 4355 64164 4359 64220
rect 4295 64160 4359 64164
rect 4375 64220 4439 64224
rect 4375 64164 4379 64220
rect 4379 64164 4435 64220
rect 4435 64164 4439 64220
rect 4375 64160 4439 64164
rect 4455 64220 4519 64224
rect 4455 64164 4459 64220
rect 4459 64164 4515 64220
rect 4515 64164 4519 64220
rect 4455 64160 4519 64164
rect 7479 64220 7543 64224
rect 7479 64164 7483 64220
rect 7483 64164 7539 64220
rect 7539 64164 7543 64220
rect 7479 64160 7543 64164
rect 7559 64220 7623 64224
rect 7559 64164 7563 64220
rect 7563 64164 7619 64220
rect 7619 64164 7623 64220
rect 7559 64160 7623 64164
rect 7639 64220 7703 64224
rect 7639 64164 7643 64220
rect 7643 64164 7699 64220
rect 7699 64164 7703 64220
rect 7639 64160 7703 64164
rect 7719 64220 7783 64224
rect 7719 64164 7723 64220
rect 7723 64164 7779 64220
rect 7779 64164 7783 64220
rect 7719 64160 7783 64164
rect 2584 63676 2648 63680
rect 2584 63620 2588 63676
rect 2588 63620 2644 63676
rect 2644 63620 2648 63676
rect 2584 63616 2648 63620
rect 2664 63676 2728 63680
rect 2664 63620 2668 63676
rect 2668 63620 2724 63676
rect 2724 63620 2728 63676
rect 2664 63616 2728 63620
rect 2744 63676 2808 63680
rect 2744 63620 2748 63676
rect 2748 63620 2804 63676
rect 2804 63620 2808 63676
rect 2744 63616 2808 63620
rect 2824 63676 2888 63680
rect 2824 63620 2828 63676
rect 2828 63620 2884 63676
rect 2884 63620 2888 63676
rect 2824 63616 2888 63620
rect 5847 63676 5911 63680
rect 5847 63620 5851 63676
rect 5851 63620 5907 63676
rect 5907 63620 5911 63676
rect 5847 63616 5911 63620
rect 5927 63676 5991 63680
rect 5927 63620 5931 63676
rect 5931 63620 5987 63676
rect 5987 63620 5991 63676
rect 5927 63616 5991 63620
rect 6007 63676 6071 63680
rect 6007 63620 6011 63676
rect 6011 63620 6067 63676
rect 6067 63620 6071 63676
rect 6007 63616 6071 63620
rect 6087 63676 6151 63680
rect 6087 63620 6091 63676
rect 6091 63620 6147 63676
rect 6147 63620 6151 63676
rect 6087 63616 6151 63620
rect 9111 63676 9175 63680
rect 9111 63620 9115 63676
rect 9115 63620 9171 63676
rect 9171 63620 9175 63676
rect 9111 63616 9175 63620
rect 9191 63676 9255 63680
rect 9191 63620 9195 63676
rect 9195 63620 9251 63676
rect 9251 63620 9255 63676
rect 9191 63616 9255 63620
rect 9271 63676 9335 63680
rect 9271 63620 9275 63676
rect 9275 63620 9331 63676
rect 9331 63620 9335 63676
rect 9271 63616 9335 63620
rect 9351 63676 9415 63680
rect 9351 63620 9355 63676
rect 9355 63620 9411 63676
rect 9411 63620 9415 63676
rect 9351 63616 9415 63620
rect 4215 63132 4279 63136
rect 4215 63076 4219 63132
rect 4219 63076 4275 63132
rect 4275 63076 4279 63132
rect 4215 63072 4279 63076
rect 4295 63132 4359 63136
rect 4295 63076 4299 63132
rect 4299 63076 4355 63132
rect 4355 63076 4359 63132
rect 4295 63072 4359 63076
rect 4375 63132 4439 63136
rect 4375 63076 4379 63132
rect 4379 63076 4435 63132
rect 4435 63076 4439 63132
rect 4375 63072 4439 63076
rect 4455 63132 4519 63136
rect 4455 63076 4459 63132
rect 4459 63076 4515 63132
rect 4515 63076 4519 63132
rect 4455 63072 4519 63076
rect 7479 63132 7543 63136
rect 7479 63076 7483 63132
rect 7483 63076 7539 63132
rect 7539 63076 7543 63132
rect 7479 63072 7543 63076
rect 7559 63132 7623 63136
rect 7559 63076 7563 63132
rect 7563 63076 7619 63132
rect 7619 63076 7623 63132
rect 7559 63072 7623 63076
rect 7639 63132 7703 63136
rect 7639 63076 7643 63132
rect 7643 63076 7699 63132
rect 7699 63076 7703 63132
rect 7639 63072 7703 63076
rect 7719 63132 7783 63136
rect 7719 63076 7723 63132
rect 7723 63076 7779 63132
rect 7779 63076 7783 63132
rect 7719 63072 7783 63076
rect 2584 62588 2648 62592
rect 2584 62532 2588 62588
rect 2588 62532 2644 62588
rect 2644 62532 2648 62588
rect 2584 62528 2648 62532
rect 2664 62588 2728 62592
rect 2664 62532 2668 62588
rect 2668 62532 2724 62588
rect 2724 62532 2728 62588
rect 2664 62528 2728 62532
rect 2744 62588 2808 62592
rect 2744 62532 2748 62588
rect 2748 62532 2804 62588
rect 2804 62532 2808 62588
rect 2744 62528 2808 62532
rect 2824 62588 2888 62592
rect 2824 62532 2828 62588
rect 2828 62532 2884 62588
rect 2884 62532 2888 62588
rect 2824 62528 2888 62532
rect 5847 62588 5911 62592
rect 5847 62532 5851 62588
rect 5851 62532 5907 62588
rect 5907 62532 5911 62588
rect 5847 62528 5911 62532
rect 5927 62588 5991 62592
rect 5927 62532 5931 62588
rect 5931 62532 5987 62588
rect 5987 62532 5991 62588
rect 5927 62528 5991 62532
rect 6007 62588 6071 62592
rect 6007 62532 6011 62588
rect 6011 62532 6067 62588
rect 6067 62532 6071 62588
rect 6007 62528 6071 62532
rect 6087 62588 6151 62592
rect 6087 62532 6091 62588
rect 6091 62532 6147 62588
rect 6147 62532 6151 62588
rect 6087 62528 6151 62532
rect 9111 62588 9175 62592
rect 9111 62532 9115 62588
rect 9115 62532 9171 62588
rect 9171 62532 9175 62588
rect 9111 62528 9175 62532
rect 9191 62588 9255 62592
rect 9191 62532 9195 62588
rect 9195 62532 9251 62588
rect 9251 62532 9255 62588
rect 9191 62528 9255 62532
rect 9271 62588 9335 62592
rect 9271 62532 9275 62588
rect 9275 62532 9331 62588
rect 9331 62532 9335 62588
rect 9271 62528 9335 62532
rect 9351 62588 9415 62592
rect 9351 62532 9355 62588
rect 9355 62532 9411 62588
rect 9411 62532 9415 62588
rect 9351 62528 9415 62532
rect 4215 62044 4279 62048
rect 4215 61988 4219 62044
rect 4219 61988 4275 62044
rect 4275 61988 4279 62044
rect 4215 61984 4279 61988
rect 4295 62044 4359 62048
rect 4295 61988 4299 62044
rect 4299 61988 4355 62044
rect 4355 61988 4359 62044
rect 4295 61984 4359 61988
rect 4375 62044 4439 62048
rect 4375 61988 4379 62044
rect 4379 61988 4435 62044
rect 4435 61988 4439 62044
rect 4375 61984 4439 61988
rect 4455 62044 4519 62048
rect 4455 61988 4459 62044
rect 4459 61988 4515 62044
rect 4515 61988 4519 62044
rect 4455 61984 4519 61988
rect 7479 62044 7543 62048
rect 7479 61988 7483 62044
rect 7483 61988 7539 62044
rect 7539 61988 7543 62044
rect 7479 61984 7543 61988
rect 7559 62044 7623 62048
rect 7559 61988 7563 62044
rect 7563 61988 7619 62044
rect 7619 61988 7623 62044
rect 7559 61984 7623 61988
rect 7639 62044 7703 62048
rect 7639 61988 7643 62044
rect 7643 61988 7699 62044
rect 7699 61988 7703 62044
rect 7639 61984 7703 61988
rect 7719 62044 7783 62048
rect 7719 61988 7723 62044
rect 7723 61988 7779 62044
rect 7779 61988 7783 62044
rect 7719 61984 7783 61988
rect 2584 61500 2648 61504
rect 2584 61444 2588 61500
rect 2588 61444 2644 61500
rect 2644 61444 2648 61500
rect 2584 61440 2648 61444
rect 2664 61500 2728 61504
rect 2664 61444 2668 61500
rect 2668 61444 2724 61500
rect 2724 61444 2728 61500
rect 2664 61440 2728 61444
rect 2744 61500 2808 61504
rect 2744 61444 2748 61500
rect 2748 61444 2804 61500
rect 2804 61444 2808 61500
rect 2744 61440 2808 61444
rect 2824 61500 2888 61504
rect 2824 61444 2828 61500
rect 2828 61444 2884 61500
rect 2884 61444 2888 61500
rect 2824 61440 2888 61444
rect 5847 61500 5911 61504
rect 5847 61444 5851 61500
rect 5851 61444 5907 61500
rect 5907 61444 5911 61500
rect 5847 61440 5911 61444
rect 5927 61500 5991 61504
rect 5927 61444 5931 61500
rect 5931 61444 5987 61500
rect 5987 61444 5991 61500
rect 5927 61440 5991 61444
rect 6007 61500 6071 61504
rect 6007 61444 6011 61500
rect 6011 61444 6067 61500
rect 6067 61444 6071 61500
rect 6007 61440 6071 61444
rect 6087 61500 6151 61504
rect 6087 61444 6091 61500
rect 6091 61444 6147 61500
rect 6147 61444 6151 61500
rect 6087 61440 6151 61444
rect 9111 61500 9175 61504
rect 9111 61444 9115 61500
rect 9115 61444 9171 61500
rect 9171 61444 9175 61500
rect 9111 61440 9175 61444
rect 9191 61500 9255 61504
rect 9191 61444 9195 61500
rect 9195 61444 9251 61500
rect 9251 61444 9255 61500
rect 9191 61440 9255 61444
rect 9271 61500 9335 61504
rect 9271 61444 9275 61500
rect 9275 61444 9331 61500
rect 9331 61444 9335 61500
rect 9271 61440 9335 61444
rect 9351 61500 9415 61504
rect 9351 61444 9355 61500
rect 9355 61444 9411 61500
rect 9411 61444 9415 61500
rect 9351 61440 9415 61444
rect 4215 60956 4279 60960
rect 4215 60900 4219 60956
rect 4219 60900 4275 60956
rect 4275 60900 4279 60956
rect 4215 60896 4279 60900
rect 4295 60956 4359 60960
rect 4295 60900 4299 60956
rect 4299 60900 4355 60956
rect 4355 60900 4359 60956
rect 4295 60896 4359 60900
rect 4375 60956 4439 60960
rect 4375 60900 4379 60956
rect 4379 60900 4435 60956
rect 4435 60900 4439 60956
rect 4375 60896 4439 60900
rect 4455 60956 4519 60960
rect 4455 60900 4459 60956
rect 4459 60900 4515 60956
rect 4515 60900 4519 60956
rect 4455 60896 4519 60900
rect 7479 60956 7543 60960
rect 7479 60900 7483 60956
rect 7483 60900 7539 60956
rect 7539 60900 7543 60956
rect 7479 60896 7543 60900
rect 7559 60956 7623 60960
rect 7559 60900 7563 60956
rect 7563 60900 7619 60956
rect 7619 60900 7623 60956
rect 7559 60896 7623 60900
rect 7639 60956 7703 60960
rect 7639 60900 7643 60956
rect 7643 60900 7699 60956
rect 7699 60900 7703 60956
rect 7639 60896 7703 60900
rect 7719 60956 7783 60960
rect 7719 60900 7723 60956
rect 7723 60900 7779 60956
rect 7779 60900 7783 60956
rect 7719 60896 7783 60900
rect 2584 60412 2648 60416
rect 2584 60356 2588 60412
rect 2588 60356 2644 60412
rect 2644 60356 2648 60412
rect 2584 60352 2648 60356
rect 2664 60412 2728 60416
rect 2664 60356 2668 60412
rect 2668 60356 2724 60412
rect 2724 60356 2728 60412
rect 2664 60352 2728 60356
rect 2744 60412 2808 60416
rect 2744 60356 2748 60412
rect 2748 60356 2804 60412
rect 2804 60356 2808 60412
rect 2744 60352 2808 60356
rect 2824 60412 2888 60416
rect 2824 60356 2828 60412
rect 2828 60356 2884 60412
rect 2884 60356 2888 60412
rect 2824 60352 2888 60356
rect 5847 60412 5911 60416
rect 5847 60356 5851 60412
rect 5851 60356 5907 60412
rect 5907 60356 5911 60412
rect 5847 60352 5911 60356
rect 5927 60412 5991 60416
rect 5927 60356 5931 60412
rect 5931 60356 5987 60412
rect 5987 60356 5991 60412
rect 5927 60352 5991 60356
rect 6007 60412 6071 60416
rect 6007 60356 6011 60412
rect 6011 60356 6067 60412
rect 6067 60356 6071 60412
rect 6007 60352 6071 60356
rect 6087 60412 6151 60416
rect 6087 60356 6091 60412
rect 6091 60356 6147 60412
rect 6147 60356 6151 60412
rect 6087 60352 6151 60356
rect 9111 60412 9175 60416
rect 9111 60356 9115 60412
rect 9115 60356 9171 60412
rect 9171 60356 9175 60412
rect 9111 60352 9175 60356
rect 9191 60412 9255 60416
rect 9191 60356 9195 60412
rect 9195 60356 9251 60412
rect 9251 60356 9255 60412
rect 9191 60352 9255 60356
rect 9271 60412 9335 60416
rect 9271 60356 9275 60412
rect 9275 60356 9331 60412
rect 9331 60356 9335 60412
rect 9271 60352 9335 60356
rect 9351 60412 9415 60416
rect 9351 60356 9355 60412
rect 9355 60356 9411 60412
rect 9411 60356 9415 60412
rect 9351 60352 9415 60356
rect 4215 59868 4279 59872
rect 4215 59812 4219 59868
rect 4219 59812 4275 59868
rect 4275 59812 4279 59868
rect 4215 59808 4279 59812
rect 4295 59868 4359 59872
rect 4295 59812 4299 59868
rect 4299 59812 4355 59868
rect 4355 59812 4359 59868
rect 4295 59808 4359 59812
rect 4375 59868 4439 59872
rect 4375 59812 4379 59868
rect 4379 59812 4435 59868
rect 4435 59812 4439 59868
rect 4375 59808 4439 59812
rect 4455 59868 4519 59872
rect 4455 59812 4459 59868
rect 4459 59812 4515 59868
rect 4515 59812 4519 59868
rect 4455 59808 4519 59812
rect 7479 59868 7543 59872
rect 7479 59812 7483 59868
rect 7483 59812 7539 59868
rect 7539 59812 7543 59868
rect 7479 59808 7543 59812
rect 7559 59868 7623 59872
rect 7559 59812 7563 59868
rect 7563 59812 7619 59868
rect 7619 59812 7623 59868
rect 7559 59808 7623 59812
rect 7639 59868 7703 59872
rect 7639 59812 7643 59868
rect 7643 59812 7699 59868
rect 7699 59812 7703 59868
rect 7639 59808 7703 59812
rect 7719 59868 7783 59872
rect 7719 59812 7723 59868
rect 7723 59812 7779 59868
rect 7779 59812 7783 59868
rect 7719 59808 7783 59812
rect 1716 59332 1780 59396
rect 2584 59324 2648 59328
rect 2584 59268 2588 59324
rect 2588 59268 2644 59324
rect 2644 59268 2648 59324
rect 2584 59264 2648 59268
rect 2664 59324 2728 59328
rect 2664 59268 2668 59324
rect 2668 59268 2724 59324
rect 2724 59268 2728 59324
rect 2664 59264 2728 59268
rect 2744 59324 2808 59328
rect 2744 59268 2748 59324
rect 2748 59268 2804 59324
rect 2804 59268 2808 59324
rect 2744 59264 2808 59268
rect 2824 59324 2888 59328
rect 2824 59268 2828 59324
rect 2828 59268 2884 59324
rect 2884 59268 2888 59324
rect 2824 59264 2888 59268
rect 5847 59324 5911 59328
rect 5847 59268 5851 59324
rect 5851 59268 5907 59324
rect 5907 59268 5911 59324
rect 5847 59264 5911 59268
rect 5927 59324 5991 59328
rect 5927 59268 5931 59324
rect 5931 59268 5987 59324
rect 5987 59268 5991 59324
rect 5927 59264 5991 59268
rect 6007 59324 6071 59328
rect 6007 59268 6011 59324
rect 6011 59268 6067 59324
rect 6067 59268 6071 59324
rect 6007 59264 6071 59268
rect 6087 59324 6151 59328
rect 6087 59268 6091 59324
rect 6091 59268 6147 59324
rect 6147 59268 6151 59324
rect 6087 59264 6151 59268
rect 9111 59324 9175 59328
rect 9111 59268 9115 59324
rect 9115 59268 9171 59324
rect 9171 59268 9175 59324
rect 9111 59264 9175 59268
rect 9191 59324 9255 59328
rect 9191 59268 9195 59324
rect 9195 59268 9251 59324
rect 9251 59268 9255 59324
rect 9191 59264 9255 59268
rect 9271 59324 9335 59328
rect 9271 59268 9275 59324
rect 9275 59268 9331 59324
rect 9331 59268 9335 59324
rect 9271 59264 9335 59268
rect 9351 59324 9415 59328
rect 9351 59268 9355 59324
rect 9355 59268 9411 59324
rect 9411 59268 9415 59324
rect 9351 59264 9415 59268
rect 4215 58780 4279 58784
rect 4215 58724 4219 58780
rect 4219 58724 4275 58780
rect 4275 58724 4279 58780
rect 4215 58720 4279 58724
rect 4295 58780 4359 58784
rect 4295 58724 4299 58780
rect 4299 58724 4355 58780
rect 4355 58724 4359 58780
rect 4295 58720 4359 58724
rect 4375 58780 4439 58784
rect 4375 58724 4379 58780
rect 4379 58724 4435 58780
rect 4435 58724 4439 58780
rect 4375 58720 4439 58724
rect 4455 58780 4519 58784
rect 4455 58724 4459 58780
rect 4459 58724 4515 58780
rect 4515 58724 4519 58780
rect 4455 58720 4519 58724
rect 7479 58780 7543 58784
rect 7479 58724 7483 58780
rect 7483 58724 7539 58780
rect 7539 58724 7543 58780
rect 7479 58720 7543 58724
rect 7559 58780 7623 58784
rect 7559 58724 7563 58780
rect 7563 58724 7619 58780
rect 7619 58724 7623 58780
rect 7559 58720 7623 58724
rect 7639 58780 7703 58784
rect 7639 58724 7643 58780
rect 7643 58724 7699 58780
rect 7699 58724 7703 58780
rect 7639 58720 7703 58724
rect 7719 58780 7783 58784
rect 7719 58724 7723 58780
rect 7723 58724 7779 58780
rect 7779 58724 7783 58780
rect 7719 58720 7783 58724
rect 2584 58236 2648 58240
rect 2584 58180 2588 58236
rect 2588 58180 2644 58236
rect 2644 58180 2648 58236
rect 2584 58176 2648 58180
rect 2664 58236 2728 58240
rect 2664 58180 2668 58236
rect 2668 58180 2724 58236
rect 2724 58180 2728 58236
rect 2664 58176 2728 58180
rect 2744 58236 2808 58240
rect 2744 58180 2748 58236
rect 2748 58180 2804 58236
rect 2804 58180 2808 58236
rect 2744 58176 2808 58180
rect 2824 58236 2888 58240
rect 2824 58180 2828 58236
rect 2828 58180 2884 58236
rect 2884 58180 2888 58236
rect 2824 58176 2888 58180
rect 5847 58236 5911 58240
rect 5847 58180 5851 58236
rect 5851 58180 5907 58236
rect 5907 58180 5911 58236
rect 5847 58176 5911 58180
rect 5927 58236 5991 58240
rect 5927 58180 5931 58236
rect 5931 58180 5987 58236
rect 5987 58180 5991 58236
rect 5927 58176 5991 58180
rect 6007 58236 6071 58240
rect 6007 58180 6011 58236
rect 6011 58180 6067 58236
rect 6067 58180 6071 58236
rect 6007 58176 6071 58180
rect 6087 58236 6151 58240
rect 6087 58180 6091 58236
rect 6091 58180 6147 58236
rect 6147 58180 6151 58236
rect 6087 58176 6151 58180
rect 9111 58236 9175 58240
rect 9111 58180 9115 58236
rect 9115 58180 9171 58236
rect 9171 58180 9175 58236
rect 9111 58176 9175 58180
rect 9191 58236 9255 58240
rect 9191 58180 9195 58236
rect 9195 58180 9251 58236
rect 9251 58180 9255 58236
rect 9191 58176 9255 58180
rect 9271 58236 9335 58240
rect 9271 58180 9275 58236
rect 9275 58180 9331 58236
rect 9331 58180 9335 58236
rect 9271 58176 9335 58180
rect 9351 58236 9415 58240
rect 9351 58180 9355 58236
rect 9355 58180 9411 58236
rect 9411 58180 9415 58236
rect 9351 58176 9415 58180
rect 4215 57692 4279 57696
rect 4215 57636 4219 57692
rect 4219 57636 4275 57692
rect 4275 57636 4279 57692
rect 4215 57632 4279 57636
rect 4295 57692 4359 57696
rect 4295 57636 4299 57692
rect 4299 57636 4355 57692
rect 4355 57636 4359 57692
rect 4295 57632 4359 57636
rect 4375 57692 4439 57696
rect 4375 57636 4379 57692
rect 4379 57636 4435 57692
rect 4435 57636 4439 57692
rect 4375 57632 4439 57636
rect 4455 57692 4519 57696
rect 4455 57636 4459 57692
rect 4459 57636 4515 57692
rect 4515 57636 4519 57692
rect 4455 57632 4519 57636
rect 7479 57692 7543 57696
rect 7479 57636 7483 57692
rect 7483 57636 7539 57692
rect 7539 57636 7543 57692
rect 7479 57632 7543 57636
rect 7559 57692 7623 57696
rect 7559 57636 7563 57692
rect 7563 57636 7619 57692
rect 7619 57636 7623 57692
rect 7559 57632 7623 57636
rect 7639 57692 7703 57696
rect 7639 57636 7643 57692
rect 7643 57636 7699 57692
rect 7699 57636 7703 57692
rect 7639 57632 7703 57636
rect 7719 57692 7783 57696
rect 7719 57636 7723 57692
rect 7723 57636 7779 57692
rect 7779 57636 7783 57692
rect 7719 57632 7783 57636
rect 2584 57148 2648 57152
rect 2584 57092 2588 57148
rect 2588 57092 2644 57148
rect 2644 57092 2648 57148
rect 2584 57088 2648 57092
rect 2664 57148 2728 57152
rect 2664 57092 2668 57148
rect 2668 57092 2724 57148
rect 2724 57092 2728 57148
rect 2664 57088 2728 57092
rect 2744 57148 2808 57152
rect 2744 57092 2748 57148
rect 2748 57092 2804 57148
rect 2804 57092 2808 57148
rect 2744 57088 2808 57092
rect 2824 57148 2888 57152
rect 2824 57092 2828 57148
rect 2828 57092 2884 57148
rect 2884 57092 2888 57148
rect 2824 57088 2888 57092
rect 5847 57148 5911 57152
rect 5847 57092 5851 57148
rect 5851 57092 5907 57148
rect 5907 57092 5911 57148
rect 5847 57088 5911 57092
rect 5927 57148 5991 57152
rect 5927 57092 5931 57148
rect 5931 57092 5987 57148
rect 5987 57092 5991 57148
rect 5927 57088 5991 57092
rect 6007 57148 6071 57152
rect 6007 57092 6011 57148
rect 6011 57092 6067 57148
rect 6067 57092 6071 57148
rect 6007 57088 6071 57092
rect 6087 57148 6151 57152
rect 6087 57092 6091 57148
rect 6091 57092 6147 57148
rect 6147 57092 6151 57148
rect 6087 57088 6151 57092
rect 9111 57148 9175 57152
rect 9111 57092 9115 57148
rect 9115 57092 9171 57148
rect 9171 57092 9175 57148
rect 9111 57088 9175 57092
rect 9191 57148 9255 57152
rect 9191 57092 9195 57148
rect 9195 57092 9251 57148
rect 9251 57092 9255 57148
rect 9191 57088 9255 57092
rect 9271 57148 9335 57152
rect 9271 57092 9275 57148
rect 9275 57092 9331 57148
rect 9331 57092 9335 57148
rect 9271 57088 9335 57092
rect 9351 57148 9415 57152
rect 9351 57092 9355 57148
rect 9355 57092 9411 57148
rect 9411 57092 9415 57148
rect 9351 57088 9415 57092
rect 4215 56604 4279 56608
rect 4215 56548 4219 56604
rect 4219 56548 4275 56604
rect 4275 56548 4279 56604
rect 4215 56544 4279 56548
rect 4295 56604 4359 56608
rect 4295 56548 4299 56604
rect 4299 56548 4355 56604
rect 4355 56548 4359 56604
rect 4295 56544 4359 56548
rect 4375 56604 4439 56608
rect 4375 56548 4379 56604
rect 4379 56548 4435 56604
rect 4435 56548 4439 56604
rect 4375 56544 4439 56548
rect 4455 56604 4519 56608
rect 4455 56548 4459 56604
rect 4459 56548 4515 56604
rect 4515 56548 4519 56604
rect 4455 56544 4519 56548
rect 7479 56604 7543 56608
rect 7479 56548 7483 56604
rect 7483 56548 7539 56604
rect 7539 56548 7543 56604
rect 7479 56544 7543 56548
rect 7559 56604 7623 56608
rect 7559 56548 7563 56604
rect 7563 56548 7619 56604
rect 7619 56548 7623 56604
rect 7559 56544 7623 56548
rect 7639 56604 7703 56608
rect 7639 56548 7643 56604
rect 7643 56548 7699 56604
rect 7699 56548 7703 56604
rect 7639 56544 7703 56548
rect 7719 56604 7783 56608
rect 7719 56548 7723 56604
rect 7723 56548 7779 56604
rect 7779 56548 7783 56604
rect 7719 56544 7783 56548
rect 2584 56060 2648 56064
rect 2584 56004 2588 56060
rect 2588 56004 2644 56060
rect 2644 56004 2648 56060
rect 2584 56000 2648 56004
rect 2664 56060 2728 56064
rect 2664 56004 2668 56060
rect 2668 56004 2724 56060
rect 2724 56004 2728 56060
rect 2664 56000 2728 56004
rect 2744 56060 2808 56064
rect 2744 56004 2748 56060
rect 2748 56004 2804 56060
rect 2804 56004 2808 56060
rect 2744 56000 2808 56004
rect 2824 56060 2888 56064
rect 2824 56004 2828 56060
rect 2828 56004 2884 56060
rect 2884 56004 2888 56060
rect 2824 56000 2888 56004
rect 5847 56060 5911 56064
rect 5847 56004 5851 56060
rect 5851 56004 5907 56060
rect 5907 56004 5911 56060
rect 5847 56000 5911 56004
rect 5927 56060 5991 56064
rect 5927 56004 5931 56060
rect 5931 56004 5987 56060
rect 5987 56004 5991 56060
rect 5927 56000 5991 56004
rect 6007 56060 6071 56064
rect 6007 56004 6011 56060
rect 6011 56004 6067 56060
rect 6067 56004 6071 56060
rect 6007 56000 6071 56004
rect 6087 56060 6151 56064
rect 6087 56004 6091 56060
rect 6091 56004 6147 56060
rect 6147 56004 6151 56060
rect 6087 56000 6151 56004
rect 9111 56060 9175 56064
rect 9111 56004 9115 56060
rect 9115 56004 9171 56060
rect 9171 56004 9175 56060
rect 9111 56000 9175 56004
rect 9191 56060 9255 56064
rect 9191 56004 9195 56060
rect 9195 56004 9251 56060
rect 9251 56004 9255 56060
rect 9191 56000 9255 56004
rect 9271 56060 9335 56064
rect 9271 56004 9275 56060
rect 9275 56004 9331 56060
rect 9331 56004 9335 56060
rect 9271 56000 9335 56004
rect 9351 56060 9415 56064
rect 9351 56004 9355 56060
rect 9355 56004 9411 56060
rect 9411 56004 9415 56060
rect 9351 56000 9415 56004
rect 4215 55516 4279 55520
rect 4215 55460 4219 55516
rect 4219 55460 4275 55516
rect 4275 55460 4279 55516
rect 4215 55456 4279 55460
rect 4295 55516 4359 55520
rect 4295 55460 4299 55516
rect 4299 55460 4355 55516
rect 4355 55460 4359 55516
rect 4295 55456 4359 55460
rect 4375 55516 4439 55520
rect 4375 55460 4379 55516
rect 4379 55460 4435 55516
rect 4435 55460 4439 55516
rect 4375 55456 4439 55460
rect 4455 55516 4519 55520
rect 4455 55460 4459 55516
rect 4459 55460 4515 55516
rect 4515 55460 4519 55516
rect 4455 55456 4519 55460
rect 7479 55516 7543 55520
rect 7479 55460 7483 55516
rect 7483 55460 7539 55516
rect 7539 55460 7543 55516
rect 7479 55456 7543 55460
rect 7559 55516 7623 55520
rect 7559 55460 7563 55516
rect 7563 55460 7619 55516
rect 7619 55460 7623 55516
rect 7559 55456 7623 55460
rect 7639 55516 7703 55520
rect 7639 55460 7643 55516
rect 7643 55460 7699 55516
rect 7699 55460 7703 55516
rect 7639 55456 7703 55460
rect 7719 55516 7783 55520
rect 7719 55460 7723 55516
rect 7723 55460 7779 55516
rect 7779 55460 7783 55516
rect 7719 55456 7783 55460
rect 2584 54972 2648 54976
rect 2584 54916 2588 54972
rect 2588 54916 2644 54972
rect 2644 54916 2648 54972
rect 2584 54912 2648 54916
rect 2664 54972 2728 54976
rect 2664 54916 2668 54972
rect 2668 54916 2724 54972
rect 2724 54916 2728 54972
rect 2664 54912 2728 54916
rect 2744 54972 2808 54976
rect 2744 54916 2748 54972
rect 2748 54916 2804 54972
rect 2804 54916 2808 54972
rect 2744 54912 2808 54916
rect 2824 54972 2888 54976
rect 2824 54916 2828 54972
rect 2828 54916 2884 54972
rect 2884 54916 2888 54972
rect 2824 54912 2888 54916
rect 5847 54972 5911 54976
rect 5847 54916 5851 54972
rect 5851 54916 5907 54972
rect 5907 54916 5911 54972
rect 5847 54912 5911 54916
rect 5927 54972 5991 54976
rect 5927 54916 5931 54972
rect 5931 54916 5987 54972
rect 5987 54916 5991 54972
rect 5927 54912 5991 54916
rect 6007 54972 6071 54976
rect 6007 54916 6011 54972
rect 6011 54916 6067 54972
rect 6067 54916 6071 54972
rect 6007 54912 6071 54916
rect 6087 54972 6151 54976
rect 6087 54916 6091 54972
rect 6091 54916 6147 54972
rect 6147 54916 6151 54972
rect 6087 54912 6151 54916
rect 9111 54972 9175 54976
rect 9111 54916 9115 54972
rect 9115 54916 9171 54972
rect 9171 54916 9175 54972
rect 9111 54912 9175 54916
rect 9191 54972 9255 54976
rect 9191 54916 9195 54972
rect 9195 54916 9251 54972
rect 9251 54916 9255 54972
rect 9191 54912 9255 54916
rect 9271 54972 9335 54976
rect 9271 54916 9275 54972
rect 9275 54916 9331 54972
rect 9331 54916 9335 54972
rect 9271 54912 9335 54916
rect 9351 54972 9415 54976
rect 9351 54916 9355 54972
rect 9355 54916 9411 54972
rect 9411 54916 9415 54972
rect 9351 54912 9415 54916
rect 4215 54428 4279 54432
rect 4215 54372 4219 54428
rect 4219 54372 4275 54428
rect 4275 54372 4279 54428
rect 4215 54368 4279 54372
rect 4295 54428 4359 54432
rect 4295 54372 4299 54428
rect 4299 54372 4355 54428
rect 4355 54372 4359 54428
rect 4295 54368 4359 54372
rect 4375 54428 4439 54432
rect 4375 54372 4379 54428
rect 4379 54372 4435 54428
rect 4435 54372 4439 54428
rect 4375 54368 4439 54372
rect 4455 54428 4519 54432
rect 4455 54372 4459 54428
rect 4459 54372 4515 54428
rect 4515 54372 4519 54428
rect 4455 54368 4519 54372
rect 7479 54428 7543 54432
rect 7479 54372 7483 54428
rect 7483 54372 7539 54428
rect 7539 54372 7543 54428
rect 7479 54368 7543 54372
rect 7559 54428 7623 54432
rect 7559 54372 7563 54428
rect 7563 54372 7619 54428
rect 7619 54372 7623 54428
rect 7559 54368 7623 54372
rect 7639 54428 7703 54432
rect 7639 54372 7643 54428
rect 7643 54372 7699 54428
rect 7699 54372 7703 54428
rect 7639 54368 7703 54372
rect 7719 54428 7783 54432
rect 7719 54372 7723 54428
rect 7723 54372 7779 54428
rect 7779 54372 7783 54428
rect 7719 54368 7783 54372
rect 2584 53884 2648 53888
rect 2584 53828 2588 53884
rect 2588 53828 2644 53884
rect 2644 53828 2648 53884
rect 2584 53824 2648 53828
rect 2664 53884 2728 53888
rect 2664 53828 2668 53884
rect 2668 53828 2724 53884
rect 2724 53828 2728 53884
rect 2664 53824 2728 53828
rect 2744 53884 2808 53888
rect 2744 53828 2748 53884
rect 2748 53828 2804 53884
rect 2804 53828 2808 53884
rect 2744 53824 2808 53828
rect 2824 53884 2888 53888
rect 2824 53828 2828 53884
rect 2828 53828 2884 53884
rect 2884 53828 2888 53884
rect 2824 53824 2888 53828
rect 5847 53884 5911 53888
rect 5847 53828 5851 53884
rect 5851 53828 5907 53884
rect 5907 53828 5911 53884
rect 5847 53824 5911 53828
rect 5927 53884 5991 53888
rect 5927 53828 5931 53884
rect 5931 53828 5987 53884
rect 5987 53828 5991 53884
rect 5927 53824 5991 53828
rect 6007 53884 6071 53888
rect 6007 53828 6011 53884
rect 6011 53828 6067 53884
rect 6067 53828 6071 53884
rect 6007 53824 6071 53828
rect 6087 53884 6151 53888
rect 6087 53828 6091 53884
rect 6091 53828 6147 53884
rect 6147 53828 6151 53884
rect 6087 53824 6151 53828
rect 9111 53884 9175 53888
rect 9111 53828 9115 53884
rect 9115 53828 9171 53884
rect 9171 53828 9175 53884
rect 9111 53824 9175 53828
rect 9191 53884 9255 53888
rect 9191 53828 9195 53884
rect 9195 53828 9251 53884
rect 9251 53828 9255 53884
rect 9191 53824 9255 53828
rect 9271 53884 9335 53888
rect 9271 53828 9275 53884
rect 9275 53828 9331 53884
rect 9331 53828 9335 53884
rect 9271 53824 9335 53828
rect 9351 53884 9415 53888
rect 9351 53828 9355 53884
rect 9355 53828 9411 53884
rect 9411 53828 9415 53884
rect 9351 53824 9415 53828
rect 4215 53340 4279 53344
rect 4215 53284 4219 53340
rect 4219 53284 4275 53340
rect 4275 53284 4279 53340
rect 4215 53280 4279 53284
rect 4295 53340 4359 53344
rect 4295 53284 4299 53340
rect 4299 53284 4355 53340
rect 4355 53284 4359 53340
rect 4295 53280 4359 53284
rect 4375 53340 4439 53344
rect 4375 53284 4379 53340
rect 4379 53284 4435 53340
rect 4435 53284 4439 53340
rect 4375 53280 4439 53284
rect 4455 53340 4519 53344
rect 4455 53284 4459 53340
rect 4459 53284 4515 53340
rect 4515 53284 4519 53340
rect 4455 53280 4519 53284
rect 7479 53340 7543 53344
rect 7479 53284 7483 53340
rect 7483 53284 7539 53340
rect 7539 53284 7543 53340
rect 7479 53280 7543 53284
rect 7559 53340 7623 53344
rect 7559 53284 7563 53340
rect 7563 53284 7619 53340
rect 7619 53284 7623 53340
rect 7559 53280 7623 53284
rect 7639 53340 7703 53344
rect 7639 53284 7643 53340
rect 7643 53284 7699 53340
rect 7699 53284 7703 53340
rect 7639 53280 7703 53284
rect 7719 53340 7783 53344
rect 7719 53284 7723 53340
rect 7723 53284 7779 53340
rect 7779 53284 7783 53340
rect 7719 53280 7783 53284
rect 2584 52796 2648 52800
rect 2584 52740 2588 52796
rect 2588 52740 2644 52796
rect 2644 52740 2648 52796
rect 2584 52736 2648 52740
rect 2664 52796 2728 52800
rect 2664 52740 2668 52796
rect 2668 52740 2724 52796
rect 2724 52740 2728 52796
rect 2664 52736 2728 52740
rect 2744 52796 2808 52800
rect 2744 52740 2748 52796
rect 2748 52740 2804 52796
rect 2804 52740 2808 52796
rect 2744 52736 2808 52740
rect 2824 52796 2888 52800
rect 2824 52740 2828 52796
rect 2828 52740 2884 52796
rect 2884 52740 2888 52796
rect 2824 52736 2888 52740
rect 5847 52796 5911 52800
rect 5847 52740 5851 52796
rect 5851 52740 5907 52796
rect 5907 52740 5911 52796
rect 5847 52736 5911 52740
rect 5927 52796 5991 52800
rect 5927 52740 5931 52796
rect 5931 52740 5987 52796
rect 5987 52740 5991 52796
rect 5927 52736 5991 52740
rect 6007 52796 6071 52800
rect 6007 52740 6011 52796
rect 6011 52740 6067 52796
rect 6067 52740 6071 52796
rect 6007 52736 6071 52740
rect 6087 52796 6151 52800
rect 6087 52740 6091 52796
rect 6091 52740 6147 52796
rect 6147 52740 6151 52796
rect 6087 52736 6151 52740
rect 9111 52796 9175 52800
rect 9111 52740 9115 52796
rect 9115 52740 9171 52796
rect 9171 52740 9175 52796
rect 9111 52736 9175 52740
rect 9191 52796 9255 52800
rect 9191 52740 9195 52796
rect 9195 52740 9251 52796
rect 9251 52740 9255 52796
rect 9191 52736 9255 52740
rect 9271 52796 9335 52800
rect 9271 52740 9275 52796
rect 9275 52740 9331 52796
rect 9331 52740 9335 52796
rect 9271 52736 9335 52740
rect 9351 52796 9415 52800
rect 9351 52740 9355 52796
rect 9355 52740 9411 52796
rect 9411 52740 9415 52796
rect 9351 52736 9415 52740
rect 4215 52252 4279 52256
rect 4215 52196 4219 52252
rect 4219 52196 4275 52252
rect 4275 52196 4279 52252
rect 4215 52192 4279 52196
rect 4295 52252 4359 52256
rect 4295 52196 4299 52252
rect 4299 52196 4355 52252
rect 4355 52196 4359 52252
rect 4295 52192 4359 52196
rect 4375 52252 4439 52256
rect 4375 52196 4379 52252
rect 4379 52196 4435 52252
rect 4435 52196 4439 52252
rect 4375 52192 4439 52196
rect 4455 52252 4519 52256
rect 4455 52196 4459 52252
rect 4459 52196 4515 52252
rect 4515 52196 4519 52252
rect 4455 52192 4519 52196
rect 7479 52252 7543 52256
rect 7479 52196 7483 52252
rect 7483 52196 7539 52252
rect 7539 52196 7543 52252
rect 7479 52192 7543 52196
rect 7559 52252 7623 52256
rect 7559 52196 7563 52252
rect 7563 52196 7619 52252
rect 7619 52196 7623 52252
rect 7559 52192 7623 52196
rect 7639 52252 7703 52256
rect 7639 52196 7643 52252
rect 7643 52196 7699 52252
rect 7699 52196 7703 52252
rect 7639 52192 7703 52196
rect 7719 52252 7783 52256
rect 7719 52196 7723 52252
rect 7723 52196 7779 52252
rect 7779 52196 7783 52252
rect 7719 52192 7783 52196
rect 2584 51708 2648 51712
rect 2584 51652 2588 51708
rect 2588 51652 2644 51708
rect 2644 51652 2648 51708
rect 2584 51648 2648 51652
rect 2664 51708 2728 51712
rect 2664 51652 2668 51708
rect 2668 51652 2724 51708
rect 2724 51652 2728 51708
rect 2664 51648 2728 51652
rect 2744 51708 2808 51712
rect 2744 51652 2748 51708
rect 2748 51652 2804 51708
rect 2804 51652 2808 51708
rect 2744 51648 2808 51652
rect 2824 51708 2888 51712
rect 2824 51652 2828 51708
rect 2828 51652 2884 51708
rect 2884 51652 2888 51708
rect 2824 51648 2888 51652
rect 5847 51708 5911 51712
rect 5847 51652 5851 51708
rect 5851 51652 5907 51708
rect 5907 51652 5911 51708
rect 5847 51648 5911 51652
rect 5927 51708 5991 51712
rect 5927 51652 5931 51708
rect 5931 51652 5987 51708
rect 5987 51652 5991 51708
rect 5927 51648 5991 51652
rect 6007 51708 6071 51712
rect 6007 51652 6011 51708
rect 6011 51652 6067 51708
rect 6067 51652 6071 51708
rect 6007 51648 6071 51652
rect 6087 51708 6151 51712
rect 6087 51652 6091 51708
rect 6091 51652 6147 51708
rect 6147 51652 6151 51708
rect 6087 51648 6151 51652
rect 9111 51708 9175 51712
rect 9111 51652 9115 51708
rect 9115 51652 9171 51708
rect 9171 51652 9175 51708
rect 9111 51648 9175 51652
rect 9191 51708 9255 51712
rect 9191 51652 9195 51708
rect 9195 51652 9251 51708
rect 9251 51652 9255 51708
rect 9191 51648 9255 51652
rect 9271 51708 9335 51712
rect 9271 51652 9275 51708
rect 9275 51652 9331 51708
rect 9331 51652 9335 51708
rect 9271 51648 9335 51652
rect 9351 51708 9415 51712
rect 9351 51652 9355 51708
rect 9355 51652 9411 51708
rect 9411 51652 9415 51708
rect 9351 51648 9415 51652
rect 4215 51164 4279 51168
rect 4215 51108 4219 51164
rect 4219 51108 4275 51164
rect 4275 51108 4279 51164
rect 4215 51104 4279 51108
rect 4295 51164 4359 51168
rect 4295 51108 4299 51164
rect 4299 51108 4355 51164
rect 4355 51108 4359 51164
rect 4295 51104 4359 51108
rect 4375 51164 4439 51168
rect 4375 51108 4379 51164
rect 4379 51108 4435 51164
rect 4435 51108 4439 51164
rect 4375 51104 4439 51108
rect 4455 51164 4519 51168
rect 4455 51108 4459 51164
rect 4459 51108 4515 51164
rect 4515 51108 4519 51164
rect 4455 51104 4519 51108
rect 7479 51164 7543 51168
rect 7479 51108 7483 51164
rect 7483 51108 7539 51164
rect 7539 51108 7543 51164
rect 7479 51104 7543 51108
rect 7559 51164 7623 51168
rect 7559 51108 7563 51164
rect 7563 51108 7619 51164
rect 7619 51108 7623 51164
rect 7559 51104 7623 51108
rect 7639 51164 7703 51168
rect 7639 51108 7643 51164
rect 7643 51108 7699 51164
rect 7699 51108 7703 51164
rect 7639 51104 7703 51108
rect 7719 51164 7783 51168
rect 7719 51108 7723 51164
rect 7723 51108 7779 51164
rect 7779 51108 7783 51164
rect 7719 51104 7783 51108
rect 1716 50960 1780 50964
rect 1716 50904 1730 50960
rect 1730 50904 1780 50960
rect 1716 50900 1780 50904
rect 2584 50620 2648 50624
rect 2584 50564 2588 50620
rect 2588 50564 2644 50620
rect 2644 50564 2648 50620
rect 2584 50560 2648 50564
rect 2664 50620 2728 50624
rect 2664 50564 2668 50620
rect 2668 50564 2724 50620
rect 2724 50564 2728 50620
rect 2664 50560 2728 50564
rect 2744 50620 2808 50624
rect 2744 50564 2748 50620
rect 2748 50564 2804 50620
rect 2804 50564 2808 50620
rect 2744 50560 2808 50564
rect 2824 50620 2888 50624
rect 2824 50564 2828 50620
rect 2828 50564 2884 50620
rect 2884 50564 2888 50620
rect 2824 50560 2888 50564
rect 5847 50620 5911 50624
rect 5847 50564 5851 50620
rect 5851 50564 5907 50620
rect 5907 50564 5911 50620
rect 5847 50560 5911 50564
rect 5927 50620 5991 50624
rect 5927 50564 5931 50620
rect 5931 50564 5987 50620
rect 5987 50564 5991 50620
rect 5927 50560 5991 50564
rect 6007 50620 6071 50624
rect 6007 50564 6011 50620
rect 6011 50564 6067 50620
rect 6067 50564 6071 50620
rect 6007 50560 6071 50564
rect 6087 50620 6151 50624
rect 6087 50564 6091 50620
rect 6091 50564 6147 50620
rect 6147 50564 6151 50620
rect 6087 50560 6151 50564
rect 9111 50620 9175 50624
rect 9111 50564 9115 50620
rect 9115 50564 9171 50620
rect 9171 50564 9175 50620
rect 9111 50560 9175 50564
rect 9191 50620 9255 50624
rect 9191 50564 9195 50620
rect 9195 50564 9251 50620
rect 9251 50564 9255 50620
rect 9191 50560 9255 50564
rect 9271 50620 9335 50624
rect 9271 50564 9275 50620
rect 9275 50564 9331 50620
rect 9331 50564 9335 50620
rect 9271 50560 9335 50564
rect 9351 50620 9415 50624
rect 9351 50564 9355 50620
rect 9355 50564 9411 50620
rect 9411 50564 9415 50620
rect 9351 50560 9415 50564
rect 4215 50076 4279 50080
rect 4215 50020 4219 50076
rect 4219 50020 4275 50076
rect 4275 50020 4279 50076
rect 4215 50016 4279 50020
rect 4295 50076 4359 50080
rect 4295 50020 4299 50076
rect 4299 50020 4355 50076
rect 4355 50020 4359 50076
rect 4295 50016 4359 50020
rect 4375 50076 4439 50080
rect 4375 50020 4379 50076
rect 4379 50020 4435 50076
rect 4435 50020 4439 50076
rect 4375 50016 4439 50020
rect 4455 50076 4519 50080
rect 4455 50020 4459 50076
rect 4459 50020 4515 50076
rect 4515 50020 4519 50076
rect 4455 50016 4519 50020
rect 7479 50076 7543 50080
rect 7479 50020 7483 50076
rect 7483 50020 7539 50076
rect 7539 50020 7543 50076
rect 7479 50016 7543 50020
rect 7559 50076 7623 50080
rect 7559 50020 7563 50076
rect 7563 50020 7619 50076
rect 7619 50020 7623 50076
rect 7559 50016 7623 50020
rect 7639 50076 7703 50080
rect 7639 50020 7643 50076
rect 7643 50020 7699 50076
rect 7699 50020 7703 50076
rect 7639 50016 7703 50020
rect 7719 50076 7783 50080
rect 7719 50020 7723 50076
rect 7723 50020 7779 50076
rect 7779 50020 7783 50076
rect 7719 50016 7783 50020
rect 2584 49532 2648 49536
rect 2584 49476 2588 49532
rect 2588 49476 2644 49532
rect 2644 49476 2648 49532
rect 2584 49472 2648 49476
rect 2664 49532 2728 49536
rect 2664 49476 2668 49532
rect 2668 49476 2724 49532
rect 2724 49476 2728 49532
rect 2664 49472 2728 49476
rect 2744 49532 2808 49536
rect 2744 49476 2748 49532
rect 2748 49476 2804 49532
rect 2804 49476 2808 49532
rect 2744 49472 2808 49476
rect 2824 49532 2888 49536
rect 2824 49476 2828 49532
rect 2828 49476 2884 49532
rect 2884 49476 2888 49532
rect 2824 49472 2888 49476
rect 5847 49532 5911 49536
rect 5847 49476 5851 49532
rect 5851 49476 5907 49532
rect 5907 49476 5911 49532
rect 5847 49472 5911 49476
rect 5927 49532 5991 49536
rect 5927 49476 5931 49532
rect 5931 49476 5987 49532
rect 5987 49476 5991 49532
rect 5927 49472 5991 49476
rect 6007 49532 6071 49536
rect 6007 49476 6011 49532
rect 6011 49476 6067 49532
rect 6067 49476 6071 49532
rect 6007 49472 6071 49476
rect 6087 49532 6151 49536
rect 6087 49476 6091 49532
rect 6091 49476 6147 49532
rect 6147 49476 6151 49532
rect 6087 49472 6151 49476
rect 9111 49532 9175 49536
rect 9111 49476 9115 49532
rect 9115 49476 9171 49532
rect 9171 49476 9175 49532
rect 9111 49472 9175 49476
rect 9191 49532 9255 49536
rect 9191 49476 9195 49532
rect 9195 49476 9251 49532
rect 9251 49476 9255 49532
rect 9191 49472 9255 49476
rect 9271 49532 9335 49536
rect 9271 49476 9275 49532
rect 9275 49476 9331 49532
rect 9331 49476 9335 49532
rect 9271 49472 9335 49476
rect 9351 49532 9415 49536
rect 9351 49476 9355 49532
rect 9355 49476 9411 49532
rect 9411 49476 9415 49532
rect 9351 49472 9415 49476
rect 4215 48988 4279 48992
rect 4215 48932 4219 48988
rect 4219 48932 4275 48988
rect 4275 48932 4279 48988
rect 4215 48928 4279 48932
rect 4295 48988 4359 48992
rect 4295 48932 4299 48988
rect 4299 48932 4355 48988
rect 4355 48932 4359 48988
rect 4295 48928 4359 48932
rect 4375 48988 4439 48992
rect 4375 48932 4379 48988
rect 4379 48932 4435 48988
rect 4435 48932 4439 48988
rect 4375 48928 4439 48932
rect 4455 48988 4519 48992
rect 4455 48932 4459 48988
rect 4459 48932 4515 48988
rect 4515 48932 4519 48988
rect 4455 48928 4519 48932
rect 7479 48988 7543 48992
rect 7479 48932 7483 48988
rect 7483 48932 7539 48988
rect 7539 48932 7543 48988
rect 7479 48928 7543 48932
rect 7559 48988 7623 48992
rect 7559 48932 7563 48988
rect 7563 48932 7619 48988
rect 7619 48932 7623 48988
rect 7559 48928 7623 48932
rect 7639 48988 7703 48992
rect 7639 48932 7643 48988
rect 7643 48932 7699 48988
rect 7699 48932 7703 48988
rect 7639 48928 7703 48932
rect 7719 48988 7783 48992
rect 7719 48932 7723 48988
rect 7723 48932 7779 48988
rect 7779 48932 7783 48988
rect 7719 48928 7783 48932
rect 2584 48444 2648 48448
rect 2584 48388 2588 48444
rect 2588 48388 2644 48444
rect 2644 48388 2648 48444
rect 2584 48384 2648 48388
rect 2664 48444 2728 48448
rect 2664 48388 2668 48444
rect 2668 48388 2724 48444
rect 2724 48388 2728 48444
rect 2664 48384 2728 48388
rect 2744 48444 2808 48448
rect 2744 48388 2748 48444
rect 2748 48388 2804 48444
rect 2804 48388 2808 48444
rect 2744 48384 2808 48388
rect 2824 48444 2888 48448
rect 2824 48388 2828 48444
rect 2828 48388 2884 48444
rect 2884 48388 2888 48444
rect 2824 48384 2888 48388
rect 5847 48444 5911 48448
rect 5847 48388 5851 48444
rect 5851 48388 5907 48444
rect 5907 48388 5911 48444
rect 5847 48384 5911 48388
rect 5927 48444 5991 48448
rect 5927 48388 5931 48444
rect 5931 48388 5987 48444
rect 5987 48388 5991 48444
rect 5927 48384 5991 48388
rect 6007 48444 6071 48448
rect 6007 48388 6011 48444
rect 6011 48388 6067 48444
rect 6067 48388 6071 48444
rect 6007 48384 6071 48388
rect 6087 48444 6151 48448
rect 6087 48388 6091 48444
rect 6091 48388 6147 48444
rect 6147 48388 6151 48444
rect 6087 48384 6151 48388
rect 9111 48444 9175 48448
rect 9111 48388 9115 48444
rect 9115 48388 9171 48444
rect 9171 48388 9175 48444
rect 9111 48384 9175 48388
rect 9191 48444 9255 48448
rect 9191 48388 9195 48444
rect 9195 48388 9251 48444
rect 9251 48388 9255 48444
rect 9191 48384 9255 48388
rect 9271 48444 9335 48448
rect 9271 48388 9275 48444
rect 9275 48388 9331 48444
rect 9331 48388 9335 48444
rect 9271 48384 9335 48388
rect 9351 48444 9415 48448
rect 9351 48388 9355 48444
rect 9355 48388 9411 48444
rect 9411 48388 9415 48444
rect 9351 48384 9415 48388
rect 4215 47900 4279 47904
rect 4215 47844 4219 47900
rect 4219 47844 4275 47900
rect 4275 47844 4279 47900
rect 4215 47840 4279 47844
rect 4295 47900 4359 47904
rect 4295 47844 4299 47900
rect 4299 47844 4355 47900
rect 4355 47844 4359 47900
rect 4295 47840 4359 47844
rect 4375 47900 4439 47904
rect 4375 47844 4379 47900
rect 4379 47844 4435 47900
rect 4435 47844 4439 47900
rect 4375 47840 4439 47844
rect 4455 47900 4519 47904
rect 4455 47844 4459 47900
rect 4459 47844 4515 47900
rect 4515 47844 4519 47900
rect 4455 47840 4519 47844
rect 7479 47900 7543 47904
rect 7479 47844 7483 47900
rect 7483 47844 7539 47900
rect 7539 47844 7543 47900
rect 7479 47840 7543 47844
rect 7559 47900 7623 47904
rect 7559 47844 7563 47900
rect 7563 47844 7619 47900
rect 7619 47844 7623 47900
rect 7559 47840 7623 47844
rect 7639 47900 7703 47904
rect 7639 47844 7643 47900
rect 7643 47844 7699 47900
rect 7699 47844 7703 47900
rect 7639 47840 7703 47844
rect 7719 47900 7783 47904
rect 7719 47844 7723 47900
rect 7723 47844 7779 47900
rect 7779 47844 7783 47900
rect 7719 47840 7783 47844
rect 2584 47356 2648 47360
rect 2584 47300 2588 47356
rect 2588 47300 2644 47356
rect 2644 47300 2648 47356
rect 2584 47296 2648 47300
rect 2664 47356 2728 47360
rect 2664 47300 2668 47356
rect 2668 47300 2724 47356
rect 2724 47300 2728 47356
rect 2664 47296 2728 47300
rect 2744 47356 2808 47360
rect 2744 47300 2748 47356
rect 2748 47300 2804 47356
rect 2804 47300 2808 47356
rect 2744 47296 2808 47300
rect 2824 47356 2888 47360
rect 2824 47300 2828 47356
rect 2828 47300 2884 47356
rect 2884 47300 2888 47356
rect 2824 47296 2888 47300
rect 5847 47356 5911 47360
rect 5847 47300 5851 47356
rect 5851 47300 5907 47356
rect 5907 47300 5911 47356
rect 5847 47296 5911 47300
rect 5927 47356 5991 47360
rect 5927 47300 5931 47356
rect 5931 47300 5987 47356
rect 5987 47300 5991 47356
rect 5927 47296 5991 47300
rect 6007 47356 6071 47360
rect 6007 47300 6011 47356
rect 6011 47300 6067 47356
rect 6067 47300 6071 47356
rect 6007 47296 6071 47300
rect 6087 47356 6151 47360
rect 6087 47300 6091 47356
rect 6091 47300 6147 47356
rect 6147 47300 6151 47356
rect 6087 47296 6151 47300
rect 9111 47356 9175 47360
rect 9111 47300 9115 47356
rect 9115 47300 9171 47356
rect 9171 47300 9175 47356
rect 9111 47296 9175 47300
rect 9191 47356 9255 47360
rect 9191 47300 9195 47356
rect 9195 47300 9251 47356
rect 9251 47300 9255 47356
rect 9191 47296 9255 47300
rect 9271 47356 9335 47360
rect 9271 47300 9275 47356
rect 9275 47300 9331 47356
rect 9331 47300 9335 47356
rect 9271 47296 9335 47300
rect 9351 47356 9415 47360
rect 9351 47300 9355 47356
rect 9355 47300 9411 47356
rect 9411 47300 9415 47356
rect 9351 47296 9415 47300
rect 3924 47152 3988 47156
rect 3924 47096 3974 47152
rect 3974 47096 3988 47152
rect 3924 47092 3988 47096
rect 4215 46812 4279 46816
rect 4215 46756 4219 46812
rect 4219 46756 4275 46812
rect 4275 46756 4279 46812
rect 4215 46752 4279 46756
rect 4295 46812 4359 46816
rect 4295 46756 4299 46812
rect 4299 46756 4355 46812
rect 4355 46756 4359 46812
rect 4295 46752 4359 46756
rect 4375 46812 4439 46816
rect 4375 46756 4379 46812
rect 4379 46756 4435 46812
rect 4435 46756 4439 46812
rect 4375 46752 4439 46756
rect 4455 46812 4519 46816
rect 4455 46756 4459 46812
rect 4459 46756 4515 46812
rect 4515 46756 4519 46812
rect 4455 46752 4519 46756
rect 7479 46812 7543 46816
rect 7479 46756 7483 46812
rect 7483 46756 7539 46812
rect 7539 46756 7543 46812
rect 7479 46752 7543 46756
rect 7559 46812 7623 46816
rect 7559 46756 7563 46812
rect 7563 46756 7619 46812
rect 7619 46756 7623 46812
rect 7559 46752 7623 46756
rect 7639 46812 7703 46816
rect 7639 46756 7643 46812
rect 7643 46756 7699 46812
rect 7699 46756 7703 46812
rect 7639 46752 7703 46756
rect 7719 46812 7783 46816
rect 7719 46756 7723 46812
rect 7723 46756 7779 46812
rect 7779 46756 7783 46812
rect 7719 46752 7783 46756
rect 2584 46268 2648 46272
rect 2584 46212 2588 46268
rect 2588 46212 2644 46268
rect 2644 46212 2648 46268
rect 2584 46208 2648 46212
rect 2664 46268 2728 46272
rect 2664 46212 2668 46268
rect 2668 46212 2724 46268
rect 2724 46212 2728 46268
rect 2664 46208 2728 46212
rect 2744 46268 2808 46272
rect 2744 46212 2748 46268
rect 2748 46212 2804 46268
rect 2804 46212 2808 46268
rect 2744 46208 2808 46212
rect 2824 46268 2888 46272
rect 2824 46212 2828 46268
rect 2828 46212 2884 46268
rect 2884 46212 2888 46268
rect 2824 46208 2888 46212
rect 5847 46268 5911 46272
rect 5847 46212 5851 46268
rect 5851 46212 5907 46268
rect 5907 46212 5911 46268
rect 5847 46208 5911 46212
rect 5927 46268 5991 46272
rect 5927 46212 5931 46268
rect 5931 46212 5987 46268
rect 5987 46212 5991 46268
rect 5927 46208 5991 46212
rect 6007 46268 6071 46272
rect 6007 46212 6011 46268
rect 6011 46212 6067 46268
rect 6067 46212 6071 46268
rect 6007 46208 6071 46212
rect 6087 46268 6151 46272
rect 6087 46212 6091 46268
rect 6091 46212 6147 46268
rect 6147 46212 6151 46268
rect 6087 46208 6151 46212
rect 9111 46268 9175 46272
rect 9111 46212 9115 46268
rect 9115 46212 9171 46268
rect 9171 46212 9175 46268
rect 9111 46208 9175 46212
rect 9191 46268 9255 46272
rect 9191 46212 9195 46268
rect 9195 46212 9251 46268
rect 9251 46212 9255 46268
rect 9191 46208 9255 46212
rect 9271 46268 9335 46272
rect 9271 46212 9275 46268
rect 9275 46212 9331 46268
rect 9331 46212 9335 46268
rect 9271 46208 9335 46212
rect 9351 46268 9415 46272
rect 9351 46212 9355 46268
rect 9355 46212 9411 46268
rect 9411 46212 9415 46268
rect 9351 46208 9415 46212
rect 4215 45724 4279 45728
rect 4215 45668 4219 45724
rect 4219 45668 4275 45724
rect 4275 45668 4279 45724
rect 4215 45664 4279 45668
rect 4295 45724 4359 45728
rect 4295 45668 4299 45724
rect 4299 45668 4355 45724
rect 4355 45668 4359 45724
rect 4295 45664 4359 45668
rect 4375 45724 4439 45728
rect 4375 45668 4379 45724
rect 4379 45668 4435 45724
rect 4435 45668 4439 45724
rect 4375 45664 4439 45668
rect 4455 45724 4519 45728
rect 4455 45668 4459 45724
rect 4459 45668 4515 45724
rect 4515 45668 4519 45724
rect 4455 45664 4519 45668
rect 7479 45724 7543 45728
rect 7479 45668 7483 45724
rect 7483 45668 7539 45724
rect 7539 45668 7543 45724
rect 7479 45664 7543 45668
rect 7559 45724 7623 45728
rect 7559 45668 7563 45724
rect 7563 45668 7619 45724
rect 7619 45668 7623 45724
rect 7559 45664 7623 45668
rect 7639 45724 7703 45728
rect 7639 45668 7643 45724
rect 7643 45668 7699 45724
rect 7699 45668 7703 45724
rect 7639 45664 7703 45668
rect 7719 45724 7783 45728
rect 7719 45668 7723 45724
rect 7723 45668 7779 45724
rect 7779 45668 7783 45724
rect 7719 45664 7783 45668
rect 2584 45180 2648 45184
rect 2584 45124 2588 45180
rect 2588 45124 2644 45180
rect 2644 45124 2648 45180
rect 2584 45120 2648 45124
rect 2664 45180 2728 45184
rect 2664 45124 2668 45180
rect 2668 45124 2724 45180
rect 2724 45124 2728 45180
rect 2664 45120 2728 45124
rect 2744 45180 2808 45184
rect 2744 45124 2748 45180
rect 2748 45124 2804 45180
rect 2804 45124 2808 45180
rect 2744 45120 2808 45124
rect 2824 45180 2888 45184
rect 2824 45124 2828 45180
rect 2828 45124 2884 45180
rect 2884 45124 2888 45180
rect 2824 45120 2888 45124
rect 5847 45180 5911 45184
rect 5847 45124 5851 45180
rect 5851 45124 5907 45180
rect 5907 45124 5911 45180
rect 5847 45120 5911 45124
rect 5927 45180 5991 45184
rect 5927 45124 5931 45180
rect 5931 45124 5987 45180
rect 5987 45124 5991 45180
rect 5927 45120 5991 45124
rect 6007 45180 6071 45184
rect 6007 45124 6011 45180
rect 6011 45124 6067 45180
rect 6067 45124 6071 45180
rect 6007 45120 6071 45124
rect 6087 45180 6151 45184
rect 6087 45124 6091 45180
rect 6091 45124 6147 45180
rect 6147 45124 6151 45180
rect 6087 45120 6151 45124
rect 9111 45180 9175 45184
rect 9111 45124 9115 45180
rect 9115 45124 9171 45180
rect 9171 45124 9175 45180
rect 9111 45120 9175 45124
rect 9191 45180 9255 45184
rect 9191 45124 9195 45180
rect 9195 45124 9251 45180
rect 9251 45124 9255 45180
rect 9191 45120 9255 45124
rect 9271 45180 9335 45184
rect 9271 45124 9275 45180
rect 9275 45124 9331 45180
rect 9331 45124 9335 45180
rect 9271 45120 9335 45124
rect 9351 45180 9415 45184
rect 9351 45124 9355 45180
rect 9355 45124 9411 45180
rect 9411 45124 9415 45180
rect 9351 45120 9415 45124
rect 3924 45112 3988 45116
rect 3924 45056 3974 45112
rect 3974 45056 3988 45112
rect 3924 45052 3988 45056
rect 4215 44636 4279 44640
rect 4215 44580 4219 44636
rect 4219 44580 4275 44636
rect 4275 44580 4279 44636
rect 4215 44576 4279 44580
rect 4295 44636 4359 44640
rect 4295 44580 4299 44636
rect 4299 44580 4355 44636
rect 4355 44580 4359 44636
rect 4295 44576 4359 44580
rect 4375 44636 4439 44640
rect 4375 44580 4379 44636
rect 4379 44580 4435 44636
rect 4435 44580 4439 44636
rect 4375 44576 4439 44580
rect 4455 44636 4519 44640
rect 4455 44580 4459 44636
rect 4459 44580 4515 44636
rect 4515 44580 4519 44636
rect 4455 44576 4519 44580
rect 7479 44636 7543 44640
rect 7479 44580 7483 44636
rect 7483 44580 7539 44636
rect 7539 44580 7543 44636
rect 7479 44576 7543 44580
rect 7559 44636 7623 44640
rect 7559 44580 7563 44636
rect 7563 44580 7619 44636
rect 7619 44580 7623 44636
rect 7559 44576 7623 44580
rect 7639 44636 7703 44640
rect 7639 44580 7643 44636
rect 7643 44580 7699 44636
rect 7699 44580 7703 44636
rect 7639 44576 7703 44580
rect 7719 44636 7783 44640
rect 7719 44580 7723 44636
rect 7723 44580 7779 44636
rect 7779 44580 7783 44636
rect 7719 44576 7783 44580
rect 2584 44092 2648 44096
rect 2584 44036 2588 44092
rect 2588 44036 2644 44092
rect 2644 44036 2648 44092
rect 2584 44032 2648 44036
rect 2664 44092 2728 44096
rect 2664 44036 2668 44092
rect 2668 44036 2724 44092
rect 2724 44036 2728 44092
rect 2664 44032 2728 44036
rect 2744 44092 2808 44096
rect 2744 44036 2748 44092
rect 2748 44036 2804 44092
rect 2804 44036 2808 44092
rect 2744 44032 2808 44036
rect 2824 44092 2888 44096
rect 2824 44036 2828 44092
rect 2828 44036 2884 44092
rect 2884 44036 2888 44092
rect 2824 44032 2888 44036
rect 5847 44092 5911 44096
rect 5847 44036 5851 44092
rect 5851 44036 5907 44092
rect 5907 44036 5911 44092
rect 5847 44032 5911 44036
rect 5927 44092 5991 44096
rect 5927 44036 5931 44092
rect 5931 44036 5987 44092
rect 5987 44036 5991 44092
rect 5927 44032 5991 44036
rect 6007 44092 6071 44096
rect 6007 44036 6011 44092
rect 6011 44036 6067 44092
rect 6067 44036 6071 44092
rect 6007 44032 6071 44036
rect 6087 44092 6151 44096
rect 6087 44036 6091 44092
rect 6091 44036 6147 44092
rect 6147 44036 6151 44092
rect 6087 44032 6151 44036
rect 9111 44092 9175 44096
rect 9111 44036 9115 44092
rect 9115 44036 9171 44092
rect 9171 44036 9175 44092
rect 9111 44032 9175 44036
rect 9191 44092 9255 44096
rect 9191 44036 9195 44092
rect 9195 44036 9251 44092
rect 9251 44036 9255 44092
rect 9191 44032 9255 44036
rect 9271 44092 9335 44096
rect 9271 44036 9275 44092
rect 9275 44036 9331 44092
rect 9331 44036 9335 44092
rect 9271 44032 9335 44036
rect 9351 44092 9415 44096
rect 9351 44036 9355 44092
rect 9355 44036 9411 44092
rect 9411 44036 9415 44092
rect 9351 44032 9415 44036
rect 4215 43548 4279 43552
rect 4215 43492 4219 43548
rect 4219 43492 4275 43548
rect 4275 43492 4279 43548
rect 4215 43488 4279 43492
rect 4295 43548 4359 43552
rect 4295 43492 4299 43548
rect 4299 43492 4355 43548
rect 4355 43492 4359 43548
rect 4295 43488 4359 43492
rect 4375 43548 4439 43552
rect 4375 43492 4379 43548
rect 4379 43492 4435 43548
rect 4435 43492 4439 43548
rect 4375 43488 4439 43492
rect 4455 43548 4519 43552
rect 4455 43492 4459 43548
rect 4459 43492 4515 43548
rect 4515 43492 4519 43548
rect 4455 43488 4519 43492
rect 7479 43548 7543 43552
rect 7479 43492 7483 43548
rect 7483 43492 7539 43548
rect 7539 43492 7543 43548
rect 7479 43488 7543 43492
rect 7559 43548 7623 43552
rect 7559 43492 7563 43548
rect 7563 43492 7619 43548
rect 7619 43492 7623 43548
rect 7559 43488 7623 43492
rect 7639 43548 7703 43552
rect 7639 43492 7643 43548
rect 7643 43492 7699 43548
rect 7699 43492 7703 43548
rect 7639 43488 7703 43492
rect 7719 43548 7783 43552
rect 7719 43492 7723 43548
rect 7723 43492 7779 43548
rect 7779 43492 7783 43548
rect 7719 43488 7783 43492
rect 2584 43004 2648 43008
rect 2584 42948 2588 43004
rect 2588 42948 2644 43004
rect 2644 42948 2648 43004
rect 2584 42944 2648 42948
rect 2664 43004 2728 43008
rect 2664 42948 2668 43004
rect 2668 42948 2724 43004
rect 2724 42948 2728 43004
rect 2664 42944 2728 42948
rect 2744 43004 2808 43008
rect 2744 42948 2748 43004
rect 2748 42948 2804 43004
rect 2804 42948 2808 43004
rect 2744 42944 2808 42948
rect 2824 43004 2888 43008
rect 2824 42948 2828 43004
rect 2828 42948 2884 43004
rect 2884 42948 2888 43004
rect 2824 42944 2888 42948
rect 5847 43004 5911 43008
rect 5847 42948 5851 43004
rect 5851 42948 5907 43004
rect 5907 42948 5911 43004
rect 5847 42944 5911 42948
rect 5927 43004 5991 43008
rect 5927 42948 5931 43004
rect 5931 42948 5987 43004
rect 5987 42948 5991 43004
rect 5927 42944 5991 42948
rect 6007 43004 6071 43008
rect 6007 42948 6011 43004
rect 6011 42948 6067 43004
rect 6067 42948 6071 43004
rect 6007 42944 6071 42948
rect 6087 43004 6151 43008
rect 6087 42948 6091 43004
rect 6091 42948 6147 43004
rect 6147 42948 6151 43004
rect 6087 42944 6151 42948
rect 9111 43004 9175 43008
rect 9111 42948 9115 43004
rect 9115 42948 9171 43004
rect 9171 42948 9175 43004
rect 9111 42944 9175 42948
rect 9191 43004 9255 43008
rect 9191 42948 9195 43004
rect 9195 42948 9251 43004
rect 9251 42948 9255 43004
rect 9191 42944 9255 42948
rect 9271 43004 9335 43008
rect 9271 42948 9275 43004
rect 9275 42948 9331 43004
rect 9331 42948 9335 43004
rect 9271 42944 9335 42948
rect 9351 43004 9415 43008
rect 9351 42948 9355 43004
rect 9355 42948 9411 43004
rect 9411 42948 9415 43004
rect 9351 42944 9415 42948
rect 4215 42460 4279 42464
rect 4215 42404 4219 42460
rect 4219 42404 4275 42460
rect 4275 42404 4279 42460
rect 4215 42400 4279 42404
rect 4295 42460 4359 42464
rect 4295 42404 4299 42460
rect 4299 42404 4355 42460
rect 4355 42404 4359 42460
rect 4295 42400 4359 42404
rect 4375 42460 4439 42464
rect 4375 42404 4379 42460
rect 4379 42404 4435 42460
rect 4435 42404 4439 42460
rect 4375 42400 4439 42404
rect 4455 42460 4519 42464
rect 4455 42404 4459 42460
rect 4459 42404 4515 42460
rect 4515 42404 4519 42460
rect 4455 42400 4519 42404
rect 7479 42460 7543 42464
rect 7479 42404 7483 42460
rect 7483 42404 7539 42460
rect 7539 42404 7543 42460
rect 7479 42400 7543 42404
rect 7559 42460 7623 42464
rect 7559 42404 7563 42460
rect 7563 42404 7619 42460
rect 7619 42404 7623 42460
rect 7559 42400 7623 42404
rect 7639 42460 7703 42464
rect 7639 42404 7643 42460
rect 7643 42404 7699 42460
rect 7699 42404 7703 42460
rect 7639 42400 7703 42404
rect 7719 42460 7783 42464
rect 7719 42404 7723 42460
rect 7723 42404 7779 42460
rect 7779 42404 7783 42460
rect 7719 42400 7783 42404
rect 2584 41916 2648 41920
rect 2584 41860 2588 41916
rect 2588 41860 2644 41916
rect 2644 41860 2648 41916
rect 2584 41856 2648 41860
rect 2664 41916 2728 41920
rect 2664 41860 2668 41916
rect 2668 41860 2724 41916
rect 2724 41860 2728 41916
rect 2664 41856 2728 41860
rect 2744 41916 2808 41920
rect 2744 41860 2748 41916
rect 2748 41860 2804 41916
rect 2804 41860 2808 41916
rect 2744 41856 2808 41860
rect 2824 41916 2888 41920
rect 2824 41860 2828 41916
rect 2828 41860 2884 41916
rect 2884 41860 2888 41916
rect 2824 41856 2888 41860
rect 5847 41916 5911 41920
rect 5847 41860 5851 41916
rect 5851 41860 5907 41916
rect 5907 41860 5911 41916
rect 5847 41856 5911 41860
rect 5927 41916 5991 41920
rect 5927 41860 5931 41916
rect 5931 41860 5987 41916
rect 5987 41860 5991 41916
rect 5927 41856 5991 41860
rect 6007 41916 6071 41920
rect 6007 41860 6011 41916
rect 6011 41860 6067 41916
rect 6067 41860 6071 41916
rect 6007 41856 6071 41860
rect 6087 41916 6151 41920
rect 6087 41860 6091 41916
rect 6091 41860 6147 41916
rect 6147 41860 6151 41916
rect 6087 41856 6151 41860
rect 9111 41916 9175 41920
rect 9111 41860 9115 41916
rect 9115 41860 9171 41916
rect 9171 41860 9175 41916
rect 9111 41856 9175 41860
rect 9191 41916 9255 41920
rect 9191 41860 9195 41916
rect 9195 41860 9251 41916
rect 9251 41860 9255 41916
rect 9191 41856 9255 41860
rect 9271 41916 9335 41920
rect 9271 41860 9275 41916
rect 9275 41860 9331 41916
rect 9331 41860 9335 41916
rect 9271 41856 9335 41860
rect 9351 41916 9415 41920
rect 9351 41860 9355 41916
rect 9355 41860 9411 41916
rect 9411 41860 9415 41916
rect 9351 41856 9415 41860
rect 3004 41788 3068 41852
rect 4660 41516 4724 41580
rect 4215 41372 4279 41376
rect 4215 41316 4219 41372
rect 4219 41316 4275 41372
rect 4275 41316 4279 41372
rect 4215 41312 4279 41316
rect 4295 41372 4359 41376
rect 4295 41316 4299 41372
rect 4299 41316 4355 41372
rect 4355 41316 4359 41372
rect 4295 41312 4359 41316
rect 4375 41372 4439 41376
rect 4375 41316 4379 41372
rect 4379 41316 4435 41372
rect 4435 41316 4439 41372
rect 4375 41312 4439 41316
rect 4455 41372 4519 41376
rect 4455 41316 4459 41372
rect 4459 41316 4515 41372
rect 4515 41316 4519 41372
rect 4455 41312 4519 41316
rect 7479 41372 7543 41376
rect 7479 41316 7483 41372
rect 7483 41316 7539 41372
rect 7539 41316 7543 41372
rect 7479 41312 7543 41316
rect 7559 41372 7623 41376
rect 7559 41316 7563 41372
rect 7563 41316 7619 41372
rect 7619 41316 7623 41372
rect 7559 41312 7623 41316
rect 7639 41372 7703 41376
rect 7639 41316 7643 41372
rect 7643 41316 7699 41372
rect 7699 41316 7703 41372
rect 7639 41312 7703 41316
rect 7719 41372 7783 41376
rect 7719 41316 7723 41372
rect 7723 41316 7779 41372
rect 7779 41316 7783 41372
rect 7719 41312 7783 41316
rect 6500 41244 6564 41308
rect 2584 40828 2648 40832
rect 2584 40772 2588 40828
rect 2588 40772 2644 40828
rect 2644 40772 2648 40828
rect 2584 40768 2648 40772
rect 2664 40828 2728 40832
rect 2664 40772 2668 40828
rect 2668 40772 2724 40828
rect 2724 40772 2728 40828
rect 2664 40768 2728 40772
rect 2744 40828 2808 40832
rect 2744 40772 2748 40828
rect 2748 40772 2804 40828
rect 2804 40772 2808 40828
rect 2744 40768 2808 40772
rect 2824 40828 2888 40832
rect 2824 40772 2828 40828
rect 2828 40772 2884 40828
rect 2884 40772 2888 40828
rect 2824 40768 2888 40772
rect 5847 40828 5911 40832
rect 5847 40772 5851 40828
rect 5851 40772 5907 40828
rect 5907 40772 5911 40828
rect 5847 40768 5911 40772
rect 5927 40828 5991 40832
rect 5927 40772 5931 40828
rect 5931 40772 5987 40828
rect 5987 40772 5991 40828
rect 5927 40768 5991 40772
rect 6007 40828 6071 40832
rect 6007 40772 6011 40828
rect 6011 40772 6067 40828
rect 6067 40772 6071 40828
rect 6007 40768 6071 40772
rect 6087 40828 6151 40832
rect 6087 40772 6091 40828
rect 6091 40772 6147 40828
rect 6147 40772 6151 40828
rect 6087 40768 6151 40772
rect 9111 40828 9175 40832
rect 9111 40772 9115 40828
rect 9115 40772 9171 40828
rect 9171 40772 9175 40828
rect 9111 40768 9175 40772
rect 9191 40828 9255 40832
rect 9191 40772 9195 40828
rect 9195 40772 9251 40828
rect 9251 40772 9255 40828
rect 9191 40768 9255 40772
rect 9271 40828 9335 40832
rect 9271 40772 9275 40828
rect 9275 40772 9331 40828
rect 9331 40772 9335 40828
rect 9271 40768 9335 40772
rect 9351 40828 9415 40832
rect 9351 40772 9355 40828
rect 9355 40772 9411 40828
rect 9411 40772 9415 40828
rect 9351 40768 9415 40772
rect 4215 40284 4279 40288
rect 4215 40228 4219 40284
rect 4219 40228 4275 40284
rect 4275 40228 4279 40284
rect 4215 40224 4279 40228
rect 4295 40284 4359 40288
rect 4295 40228 4299 40284
rect 4299 40228 4355 40284
rect 4355 40228 4359 40284
rect 4295 40224 4359 40228
rect 4375 40284 4439 40288
rect 4375 40228 4379 40284
rect 4379 40228 4435 40284
rect 4435 40228 4439 40284
rect 4375 40224 4439 40228
rect 4455 40284 4519 40288
rect 4455 40228 4459 40284
rect 4459 40228 4515 40284
rect 4515 40228 4519 40284
rect 4455 40224 4519 40228
rect 7479 40284 7543 40288
rect 7479 40228 7483 40284
rect 7483 40228 7539 40284
rect 7539 40228 7543 40284
rect 7479 40224 7543 40228
rect 7559 40284 7623 40288
rect 7559 40228 7563 40284
rect 7563 40228 7619 40284
rect 7619 40228 7623 40284
rect 7559 40224 7623 40228
rect 7639 40284 7703 40288
rect 7639 40228 7643 40284
rect 7643 40228 7699 40284
rect 7699 40228 7703 40284
rect 7639 40224 7703 40228
rect 7719 40284 7783 40288
rect 7719 40228 7723 40284
rect 7723 40228 7779 40284
rect 7779 40228 7783 40284
rect 7719 40224 7783 40228
rect 3004 40080 3068 40084
rect 3004 40024 3054 40080
rect 3054 40024 3068 40080
rect 3004 40020 3068 40024
rect 2584 39740 2648 39744
rect 2584 39684 2588 39740
rect 2588 39684 2644 39740
rect 2644 39684 2648 39740
rect 2584 39680 2648 39684
rect 2664 39740 2728 39744
rect 2664 39684 2668 39740
rect 2668 39684 2724 39740
rect 2724 39684 2728 39740
rect 2664 39680 2728 39684
rect 2744 39740 2808 39744
rect 2744 39684 2748 39740
rect 2748 39684 2804 39740
rect 2804 39684 2808 39740
rect 2744 39680 2808 39684
rect 2824 39740 2888 39744
rect 2824 39684 2828 39740
rect 2828 39684 2884 39740
rect 2884 39684 2888 39740
rect 2824 39680 2888 39684
rect 5847 39740 5911 39744
rect 5847 39684 5851 39740
rect 5851 39684 5907 39740
rect 5907 39684 5911 39740
rect 5847 39680 5911 39684
rect 5927 39740 5991 39744
rect 5927 39684 5931 39740
rect 5931 39684 5987 39740
rect 5987 39684 5991 39740
rect 5927 39680 5991 39684
rect 6007 39740 6071 39744
rect 6007 39684 6011 39740
rect 6011 39684 6067 39740
rect 6067 39684 6071 39740
rect 6007 39680 6071 39684
rect 6087 39740 6151 39744
rect 6087 39684 6091 39740
rect 6091 39684 6147 39740
rect 6147 39684 6151 39740
rect 6087 39680 6151 39684
rect 9111 39740 9175 39744
rect 9111 39684 9115 39740
rect 9115 39684 9171 39740
rect 9171 39684 9175 39740
rect 9111 39680 9175 39684
rect 9191 39740 9255 39744
rect 9191 39684 9195 39740
rect 9195 39684 9251 39740
rect 9251 39684 9255 39740
rect 9191 39680 9255 39684
rect 9271 39740 9335 39744
rect 9271 39684 9275 39740
rect 9275 39684 9331 39740
rect 9331 39684 9335 39740
rect 9271 39680 9335 39684
rect 9351 39740 9415 39744
rect 9351 39684 9355 39740
rect 9355 39684 9411 39740
rect 9411 39684 9415 39740
rect 9351 39680 9415 39684
rect 4215 39196 4279 39200
rect 4215 39140 4219 39196
rect 4219 39140 4275 39196
rect 4275 39140 4279 39196
rect 4215 39136 4279 39140
rect 4295 39196 4359 39200
rect 4295 39140 4299 39196
rect 4299 39140 4355 39196
rect 4355 39140 4359 39196
rect 4295 39136 4359 39140
rect 4375 39196 4439 39200
rect 4375 39140 4379 39196
rect 4379 39140 4435 39196
rect 4435 39140 4439 39196
rect 4375 39136 4439 39140
rect 4455 39196 4519 39200
rect 4455 39140 4459 39196
rect 4459 39140 4515 39196
rect 4515 39140 4519 39196
rect 4455 39136 4519 39140
rect 7479 39196 7543 39200
rect 7479 39140 7483 39196
rect 7483 39140 7539 39196
rect 7539 39140 7543 39196
rect 7479 39136 7543 39140
rect 7559 39196 7623 39200
rect 7559 39140 7563 39196
rect 7563 39140 7619 39196
rect 7619 39140 7623 39196
rect 7559 39136 7623 39140
rect 7639 39196 7703 39200
rect 7639 39140 7643 39196
rect 7643 39140 7699 39196
rect 7699 39140 7703 39196
rect 7639 39136 7703 39140
rect 7719 39196 7783 39200
rect 7719 39140 7723 39196
rect 7723 39140 7779 39196
rect 7779 39140 7783 39196
rect 7719 39136 7783 39140
rect 2584 38652 2648 38656
rect 2584 38596 2588 38652
rect 2588 38596 2644 38652
rect 2644 38596 2648 38652
rect 2584 38592 2648 38596
rect 2664 38652 2728 38656
rect 2664 38596 2668 38652
rect 2668 38596 2724 38652
rect 2724 38596 2728 38652
rect 2664 38592 2728 38596
rect 2744 38652 2808 38656
rect 2744 38596 2748 38652
rect 2748 38596 2804 38652
rect 2804 38596 2808 38652
rect 2744 38592 2808 38596
rect 2824 38652 2888 38656
rect 2824 38596 2828 38652
rect 2828 38596 2884 38652
rect 2884 38596 2888 38652
rect 2824 38592 2888 38596
rect 5847 38652 5911 38656
rect 5847 38596 5851 38652
rect 5851 38596 5907 38652
rect 5907 38596 5911 38652
rect 5847 38592 5911 38596
rect 5927 38652 5991 38656
rect 5927 38596 5931 38652
rect 5931 38596 5987 38652
rect 5987 38596 5991 38652
rect 5927 38592 5991 38596
rect 6007 38652 6071 38656
rect 6007 38596 6011 38652
rect 6011 38596 6067 38652
rect 6067 38596 6071 38652
rect 6007 38592 6071 38596
rect 6087 38652 6151 38656
rect 6087 38596 6091 38652
rect 6091 38596 6147 38652
rect 6147 38596 6151 38652
rect 6087 38592 6151 38596
rect 9111 38652 9175 38656
rect 9111 38596 9115 38652
rect 9115 38596 9171 38652
rect 9171 38596 9175 38652
rect 9111 38592 9175 38596
rect 9191 38652 9255 38656
rect 9191 38596 9195 38652
rect 9195 38596 9251 38652
rect 9251 38596 9255 38652
rect 9191 38592 9255 38596
rect 9271 38652 9335 38656
rect 9271 38596 9275 38652
rect 9275 38596 9331 38652
rect 9331 38596 9335 38652
rect 9271 38592 9335 38596
rect 9351 38652 9415 38656
rect 9351 38596 9355 38652
rect 9355 38596 9411 38652
rect 9411 38596 9415 38652
rect 9351 38592 9415 38596
rect 4215 38108 4279 38112
rect 4215 38052 4219 38108
rect 4219 38052 4275 38108
rect 4275 38052 4279 38108
rect 4215 38048 4279 38052
rect 4295 38108 4359 38112
rect 4295 38052 4299 38108
rect 4299 38052 4355 38108
rect 4355 38052 4359 38108
rect 4295 38048 4359 38052
rect 4375 38108 4439 38112
rect 4375 38052 4379 38108
rect 4379 38052 4435 38108
rect 4435 38052 4439 38108
rect 4375 38048 4439 38052
rect 4455 38108 4519 38112
rect 4455 38052 4459 38108
rect 4459 38052 4515 38108
rect 4515 38052 4519 38108
rect 4455 38048 4519 38052
rect 7479 38108 7543 38112
rect 7479 38052 7483 38108
rect 7483 38052 7539 38108
rect 7539 38052 7543 38108
rect 7479 38048 7543 38052
rect 7559 38108 7623 38112
rect 7559 38052 7563 38108
rect 7563 38052 7619 38108
rect 7619 38052 7623 38108
rect 7559 38048 7623 38052
rect 7639 38108 7703 38112
rect 7639 38052 7643 38108
rect 7643 38052 7699 38108
rect 7699 38052 7703 38108
rect 7639 38048 7703 38052
rect 7719 38108 7783 38112
rect 7719 38052 7723 38108
rect 7723 38052 7779 38108
rect 7779 38052 7783 38108
rect 7719 38048 7783 38052
rect 2584 37564 2648 37568
rect 2584 37508 2588 37564
rect 2588 37508 2644 37564
rect 2644 37508 2648 37564
rect 2584 37504 2648 37508
rect 2664 37564 2728 37568
rect 2664 37508 2668 37564
rect 2668 37508 2724 37564
rect 2724 37508 2728 37564
rect 2664 37504 2728 37508
rect 2744 37564 2808 37568
rect 2744 37508 2748 37564
rect 2748 37508 2804 37564
rect 2804 37508 2808 37564
rect 2744 37504 2808 37508
rect 2824 37564 2888 37568
rect 2824 37508 2828 37564
rect 2828 37508 2884 37564
rect 2884 37508 2888 37564
rect 2824 37504 2888 37508
rect 5847 37564 5911 37568
rect 5847 37508 5851 37564
rect 5851 37508 5907 37564
rect 5907 37508 5911 37564
rect 5847 37504 5911 37508
rect 5927 37564 5991 37568
rect 5927 37508 5931 37564
rect 5931 37508 5987 37564
rect 5987 37508 5991 37564
rect 5927 37504 5991 37508
rect 6007 37564 6071 37568
rect 6007 37508 6011 37564
rect 6011 37508 6067 37564
rect 6067 37508 6071 37564
rect 6007 37504 6071 37508
rect 6087 37564 6151 37568
rect 6087 37508 6091 37564
rect 6091 37508 6147 37564
rect 6147 37508 6151 37564
rect 6087 37504 6151 37508
rect 9111 37564 9175 37568
rect 9111 37508 9115 37564
rect 9115 37508 9171 37564
rect 9171 37508 9175 37564
rect 9111 37504 9175 37508
rect 9191 37564 9255 37568
rect 9191 37508 9195 37564
rect 9195 37508 9251 37564
rect 9251 37508 9255 37564
rect 9191 37504 9255 37508
rect 9271 37564 9335 37568
rect 9271 37508 9275 37564
rect 9275 37508 9331 37564
rect 9331 37508 9335 37564
rect 9271 37504 9335 37508
rect 9351 37564 9415 37568
rect 9351 37508 9355 37564
rect 9355 37508 9411 37564
rect 9411 37508 9415 37564
rect 9351 37504 9415 37508
rect 4215 37020 4279 37024
rect 4215 36964 4219 37020
rect 4219 36964 4275 37020
rect 4275 36964 4279 37020
rect 4215 36960 4279 36964
rect 4295 37020 4359 37024
rect 4295 36964 4299 37020
rect 4299 36964 4355 37020
rect 4355 36964 4359 37020
rect 4295 36960 4359 36964
rect 4375 37020 4439 37024
rect 4375 36964 4379 37020
rect 4379 36964 4435 37020
rect 4435 36964 4439 37020
rect 4375 36960 4439 36964
rect 4455 37020 4519 37024
rect 4455 36964 4459 37020
rect 4459 36964 4515 37020
rect 4515 36964 4519 37020
rect 4455 36960 4519 36964
rect 7479 37020 7543 37024
rect 7479 36964 7483 37020
rect 7483 36964 7539 37020
rect 7539 36964 7543 37020
rect 7479 36960 7543 36964
rect 7559 37020 7623 37024
rect 7559 36964 7563 37020
rect 7563 36964 7619 37020
rect 7619 36964 7623 37020
rect 7559 36960 7623 36964
rect 7639 37020 7703 37024
rect 7639 36964 7643 37020
rect 7643 36964 7699 37020
rect 7699 36964 7703 37020
rect 7639 36960 7703 36964
rect 7719 37020 7783 37024
rect 7719 36964 7723 37020
rect 7723 36964 7779 37020
rect 7779 36964 7783 37020
rect 7719 36960 7783 36964
rect 6500 36952 6564 36956
rect 6500 36896 6514 36952
rect 6514 36896 6564 36952
rect 6500 36892 6564 36896
rect 2584 36476 2648 36480
rect 2584 36420 2588 36476
rect 2588 36420 2644 36476
rect 2644 36420 2648 36476
rect 2584 36416 2648 36420
rect 2664 36476 2728 36480
rect 2664 36420 2668 36476
rect 2668 36420 2724 36476
rect 2724 36420 2728 36476
rect 2664 36416 2728 36420
rect 2744 36476 2808 36480
rect 2744 36420 2748 36476
rect 2748 36420 2804 36476
rect 2804 36420 2808 36476
rect 2744 36416 2808 36420
rect 2824 36476 2888 36480
rect 2824 36420 2828 36476
rect 2828 36420 2884 36476
rect 2884 36420 2888 36476
rect 2824 36416 2888 36420
rect 5847 36476 5911 36480
rect 5847 36420 5851 36476
rect 5851 36420 5907 36476
rect 5907 36420 5911 36476
rect 5847 36416 5911 36420
rect 5927 36476 5991 36480
rect 5927 36420 5931 36476
rect 5931 36420 5987 36476
rect 5987 36420 5991 36476
rect 5927 36416 5991 36420
rect 6007 36476 6071 36480
rect 6007 36420 6011 36476
rect 6011 36420 6067 36476
rect 6067 36420 6071 36476
rect 6007 36416 6071 36420
rect 6087 36476 6151 36480
rect 6087 36420 6091 36476
rect 6091 36420 6147 36476
rect 6147 36420 6151 36476
rect 6087 36416 6151 36420
rect 9111 36476 9175 36480
rect 9111 36420 9115 36476
rect 9115 36420 9171 36476
rect 9171 36420 9175 36476
rect 9111 36416 9175 36420
rect 9191 36476 9255 36480
rect 9191 36420 9195 36476
rect 9195 36420 9251 36476
rect 9251 36420 9255 36476
rect 9191 36416 9255 36420
rect 9271 36476 9335 36480
rect 9271 36420 9275 36476
rect 9275 36420 9331 36476
rect 9331 36420 9335 36476
rect 9271 36416 9335 36420
rect 9351 36476 9415 36480
rect 9351 36420 9355 36476
rect 9355 36420 9411 36476
rect 9411 36420 9415 36476
rect 9351 36416 9415 36420
rect 4215 35932 4279 35936
rect 4215 35876 4219 35932
rect 4219 35876 4275 35932
rect 4275 35876 4279 35932
rect 4215 35872 4279 35876
rect 4295 35932 4359 35936
rect 4295 35876 4299 35932
rect 4299 35876 4355 35932
rect 4355 35876 4359 35932
rect 4295 35872 4359 35876
rect 4375 35932 4439 35936
rect 4375 35876 4379 35932
rect 4379 35876 4435 35932
rect 4435 35876 4439 35932
rect 4375 35872 4439 35876
rect 4455 35932 4519 35936
rect 4455 35876 4459 35932
rect 4459 35876 4515 35932
rect 4515 35876 4519 35932
rect 4455 35872 4519 35876
rect 7479 35932 7543 35936
rect 7479 35876 7483 35932
rect 7483 35876 7539 35932
rect 7539 35876 7543 35932
rect 7479 35872 7543 35876
rect 7559 35932 7623 35936
rect 7559 35876 7563 35932
rect 7563 35876 7619 35932
rect 7619 35876 7623 35932
rect 7559 35872 7623 35876
rect 7639 35932 7703 35936
rect 7639 35876 7643 35932
rect 7643 35876 7699 35932
rect 7699 35876 7703 35932
rect 7639 35872 7703 35876
rect 7719 35932 7783 35936
rect 7719 35876 7723 35932
rect 7723 35876 7779 35932
rect 7779 35876 7783 35932
rect 7719 35872 7783 35876
rect 2584 35388 2648 35392
rect 2584 35332 2588 35388
rect 2588 35332 2644 35388
rect 2644 35332 2648 35388
rect 2584 35328 2648 35332
rect 2664 35388 2728 35392
rect 2664 35332 2668 35388
rect 2668 35332 2724 35388
rect 2724 35332 2728 35388
rect 2664 35328 2728 35332
rect 2744 35388 2808 35392
rect 2744 35332 2748 35388
rect 2748 35332 2804 35388
rect 2804 35332 2808 35388
rect 2744 35328 2808 35332
rect 2824 35388 2888 35392
rect 2824 35332 2828 35388
rect 2828 35332 2884 35388
rect 2884 35332 2888 35388
rect 2824 35328 2888 35332
rect 5847 35388 5911 35392
rect 5847 35332 5851 35388
rect 5851 35332 5907 35388
rect 5907 35332 5911 35388
rect 5847 35328 5911 35332
rect 5927 35388 5991 35392
rect 5927 35332 5931 35388
rect 5931 35332 5987 35388
rect 5987 35332 5991 35388
rect 5927 35328 5991 35332
rect 6007 35388 6071 35392
rect 6007 35332 6011 35388
rect 6011 35332 6067 35388
rect 6067 35332 6071 35388
rect 6007 35328 6071 35332
rect 6087 35388 6151 35392
rect 6087 35332 6091 35388
rect 6091 35332 6147 35388
rect 6147 35332 6151 35388
rect 6087 35328 6151 35332
rect 9111 35388 9175 35392
rect 9111 35332 9115 35388
rect 9115 35332 9171 35388
rect 9171 35332 9175 35388
rect 9111 35328 9175 35332
rect 9191 35388 9255 35392
rect 9191 35332 9195 35388
rect 9195 35332 9251 35388
rect 9251 35332 9255 35388
rect 9191 35328 9255 35332
rect 9271 35388 9335 35392
rect 9271 35332 9275 35388
rect 9275 35332 9331 35388
rect 9331 35332 9335 35388
rect 9271 35328 9335 35332
rect 9351 35388 9415 35392
rect 9351 35332 9355 35388
rect 9355 35332 9411 35388
rect 9411 35332 9415 35388
rect 9351 35328 9415 35332
rect 4215 34844 4279 34848
rect 4215 34788 4219 34844
rect 4219 34788 4275 34844
rect 4275 34788 4279 34844
rect 4215 34784 4279 34788
rect 4295 34844 4359 34848
rect 4295 34788 4299 34844
rect 4299 34788 4355 34844
rect 4355 34788 4359 34844
rect 4295 34784 4359 34788
rect 4375 34844 4439 34848
rect 4375 34788 4379 34844
rect 4379 34788 4435 34844
rect 4435 34788 4439 34844
rect 4375 34784 4439 34788
rect 4455 34844 4519 34848
rect 4455 34788 4459 34844
rect 4459 34788 4515 34844
rect 4515 34788 4519 34844
rect 4455 34784 4519 34788
rect 7479 34844 7543 34848
rect 7479 34788 7483 34844
rect 7483 34788 7539 34844
rect 7539 34788 7543 34844
rect 7479 34784 7543 34788
rect 7559 34844 7623 34848
rect 7559 34788 7563 34844
rect 7563 34788 7619 34844
rect 7619 34788 7623 34844
rect 7559 34784 7623 34788
rect 7639 34844 7703 34848
rect 7639 34788 7643 34844
rect 7643 34788 7699 34844
rect 7699 34788 7703 34844
rect 7639 34784 7703 34788
rect 7719 34844 7783 34848
rect 7719 34788 7723 34844
rect 7723 34788 7779 34844
rect 7779 34788 7783 34844
rect 7719 34784 7783 34788
rect 4660 34368 4724 34372
rect 4660 34312 4674 34368
rect 4674 34312 4724 34368
rect 4660 34308 4724 34312
rect 2584 34300 2648 34304
rect 2584 34244 2588 34300
rect 2588 34244 2644 34300
rect 2644 34244 2648 34300
rect 2584 34240 2648 34244
rect 2664 34300 2728 34304
rect 2664 34244 2668 34300
rect 2668 34244 2724 34300
rect 2724 34244 2728 34300
rect 2664 34240 2728 34244
rect 2744 34300 2808 34304
rect 2744 34244 2748 34300
rect 2748 34244 2804 34300
rect 2804 34244 2808 34300
rect 2744 34240 2808 34244
rect 2824 34300 2888 34304
rect 2824 34244 2828 34300
rect 2828 34244 2884 34300
rect 2884 34244 2888 34300
rect 2824 34240 2888 34244
rect 5847 34300 5911 34304
rect 5847 34244 5851 34300
rect 5851 34244 5907 34300
rect 5907 34244 5911 34300
rect 5847 34240 5911 34244
rect 5927 34300 5991 34304
rect 5927 34244 5931 34300
rect 5931 34244 5987 34300
rect 5987 34244 5991 34300
rect 5927 34240 5991 34244
rect 6007 34300 6071 34304
rect 6007 34244 6011 34300
rect 6011 34244 6067 34300
rect 6067 34244 6071 34300
rect 6007 34240 6071 34244
rect 6087 34300 6151 34304
rect 6087 34244 6091 34300
rect 6091 34244 6147 34300
rect 6147 34244 6151 34300
rect 6087 34240 6151 34244
rect 9111 34300 9175 34304
rect 9111 34244 9115 34300
rect 9115 34244 9171 34300
rect 9171 34244 9175 34300
rect 9111 34240 9175 34244
rect 9191 34300 9255 34304
rect 9191 34244 9195 34300
rect 9195 34244 9251 34300
rect 9251 34244 9255 34300
rect 9191 34240 9255 34244
rect 9271 34300 9335 34304
rect 9271 34244 9275 34300
rect 9275 34244 9331 34300
rect 9331 34244 9335 34300
rect 9271 34240 9335 34244
rect 9351 34300 9415 34304
rect 9351 34244 9355 34300
rect 9355 34244 9411 34300
rect 9411 34244 9415 34300
rect 9351 34240 9415 34244
rect 4215 33756 4279 33760
rect 4215 33700 4219 33756
rect 4219 33700 4275 33756
rect 4275 33700 4279 33756
rect 4215 33696 4279 33700
rect 4295 33756 4359 33760
rect 4295 33700 4299 33756
rect 4299 33700 4355 33756
rect 4355 33700 4359 33756
rect 4295 33696 4359 33700
rect 4375 33756 4439 33760
rect 4375 33700 4379 33756
rect 4379 33700 4435 33756
rect 4435 33700 4439 33756
rect 4375 33696 4439 33700
rect 4455 33756 4519 33760
rect 4455 33700 4459 33756
rect 4459 33700 4515 33756
rect 4515 33700 4519 33756
rect 4455 33696 4519 33700
rect 7479 33756 7543 33760
rect 7479 33700 7483 33756
rect 7483 33700 7539 33756
rect 7539 33700 7543 33756
rect 7479 33696 7543 33700
rect 7559 33756 7623 33760
rect 7559 33700 7563 33756
rect 7563 33700 7619 33756
rect 7619 33700 7623 33756
rect 7559 33696 7623 33700
rect 7639 33756 7703 33760
rect 7639 33700 7643 33756
rect 7643 33700 7699 33756
rect 7699 33700 7703 33756
rect 7639 33696 7703 33700
rect 7719 33756 7783 33760
rect 7719 33700 7723 33756
rect 7723 33700 7779 33756
rect 7779 33700 7783 33756
rect 7719 33696 7783 33700
rect 2584 33212 2648 33216
rect 2584 33156 2588 33212
rect 2588 33156 2644 33212
rect 2644 33156 2648 33212
rect 2584 33152 2648 33156
rect 2664 33212 2728 33216
rect 2664 33156 2668 33212
rect 2668 33156 2724 33212
rect 2724 33156 2728 33212
rect 2664 33152 2728 33156
rect 2744 33212 2808 33216
rect 2744 33156 2748 33212
rect 2748 33156 2804 33212
rect 2804 33156 2808 33212
rect 2744 33152 2808 33156
rect 2824 33212 2888 33216
rect 2824 33156 2828 33212
rect 2828 33156 2884 33212
rect 2884 33156 2888 33212
rect 2824 33152 2888 33156
rect 5847 33212 5911 33216
rect 5847 33156 5851 33212
rect 5851 33156 5907 33212
rect 5907 33156 5911 33212
rect 5847 33152 5911 33156
rect 5927 33212 5991 33216
rect 5927 33156 5931 33212
rect 5931 33156 5987 33212
rect 5987 33156 5991 33212
rect 5927 33152 5991 33156
rect 6007 33212 6071 33216
rect 6007 33156 6011 33212
rect 6011 33156 6067 33212
rect 6067 33156 6071 33212
rect 6007 33152 6071 33156
rect 6087 33212 6151 33216
rect 6087 33156 6091 33212
rect 6091 33156 6147 33212
rect 6147 33156 6151 33212
rect 6087 33152 6151 33156
rect 9111 33212 9175 33216
rect 9111 33156 9115 33212
rect 9115 33156 9171 33212
rect 9171 33156 9175 33212
rect 9111 33152 9175 33156
rect 9191 33212 9255 33216
rect 9191 33156 9195 33212
rect 9195 33156 9251 33212
rect 9251 33156 9255 33212
rect 9191 33152 9255 33156
rect 9271 33212 9335 33216
rect 9271 33156 9275 33212
rect 9275 33156 9331 33212
rect 9331 33156 9335 33212
rect 9271 33152 9335 33156
rect 9351 33212 9415 33216
rect 9351 33156 9355 33212
rect 9355 33156 9411 33212
rect 9411 33156 9415 33212
rect 9351 33152 9415 33156
rect 4215 32668 4279 32672
rect 4215 32612 4219 32668
rect 4219 32612 4275 32668
rect 4275 32612 4279 32668
rect 4215 32608 4279 32612
rect 4295 32668 4359 32672
rect 4295 32612 4299 32668
rect 4299 32612 4355 32668
rect 4355 32612 4359 32668
rect 4295 32608 4359 32612
rect 4375 32668 4439 32672
rect 4375 32612 4379 32668
rect 4379 32612 4435 32668
rect 4435 32612 4439 32668
rect 4375 32608 4439 32612
rect 4455 32668 4519 32672
rect 4455 32612 4459 32668
rect 4459 32612 4515 32668
rect 4515 32612 4519 32668
rect 4455 32608 4519 32612
rect 7479 32668 7543 32672
rect 7479 32612 7483 32668
rect 7483 32612 7539 32668
rect 7539 32612 7543 32668
rect 7479 32608 7543 32612
rect 7559 32668 7623 32672
rect 7559 32612 7563 32668
rect 7563 32612 7619 32668
rect 7619 32612 7623 32668
rect 7559 32608 7623 32612
rect 7639 32668 7703 32672
rect 7639 32612 7643 32668
rect 7643 32612 7699 32668
rect 7699 32612 7703 32668
rect 7639 32608 7703 32612
rect 7719 32668 7783 32672
rect 7719 32612 7723 32668
rect 7723 32612 7779 32668
rect 7779 32612 7783 32668
rect 7719 32608 7783 32612
rect 2584 32124 2648 32128
rect 2584 32068 2588 32124
rect 2588 32068 2644 32124
rect 2644 32068 2648 32124
rect 2584 32064 2648 32068
rect 2664 32124 2728 32128
rect 2664 32068 2668 32124
rect 2668 32068 2724 32124
rect 2724 32068 2728 32124
rect 2664 32064 2728 32068
rect 2744 32124 2808 32128
rect 2744 32068 2748 32124
rect 2748 32068 2804 32124
rect 2804 32068 2808 32124
rect 2744 32064 2808 32068
rect 2824 32124 2888 32128
rect 2824 32068 2828 32124
rect 2828 32068 2884 32124
rect 2884 32068 2888 32124
rect 2824 32064 2888 32068
rect 5847 32124 5911 32128
rect 5847 32068 5851 32124
rect 5851 32068 5907 32124
rect 5907 32068 5911 32124
rect 5847 32064 5911 32068
rect 5927 32124 5991 32128
rect 5927 32068 5931 32124
rect 5931 32068 5987 32124
rect 5987 32068 5991 32124
rect 5927 32064 5991 32068
rect 6007 32124 6071 32128
rect 6007 32068 6011 32124
rect 6011 32068 6067 32124
rect 6067 32068 6071 32124
rect 6007 32064 6071 32068
rect 6087 32124 6151 32128
rect 6087 32068 6091 32124
rect 6091 32068 6147 32124
rect 6147 32068 6151 32124
rect 6087 32064 6151 32068
rect 9111 32124 9175 32128
rect 9111 32068 9115 32124
rect 9115 32068 9171 32124
rect 9171 32068 9175 32124
rect 9111 32064 9175 32068
rect 9191 32124 9255 32128
rect 9191 32068 9195 32124
rect 9195 32068 9251 32124
rect 9251 32068 9255 32124
rect 9191 32064 9255 32068
rect 9271 32124 9335 32128
rect 9271 32068 9275 32124
rect 9275 32068 9331 32124
rect 9331 32068 9335 32124
rect 9271 32064 9335 32068
rect 9351 32124 9415 32128
rect 9351 32068 9355 32124
rect 9355 32068 9411 32124
rect 9411 32068 9415 32124
rect 9351 32064 9415 32068
rect 4215 31580 4279 31584
rect 4215 31524 4219 31580
rect 4219 31524 4275 31580
rect 4275 31524 4279 31580
rect 4215 31520 4279 31524
rect 4295 31580 4359 31584
rect 4295 31524 4299 31580
rect 4299 31524 4355 31580
rect 4355 31524 4359 31580
rect 4295 31520 4359 31524
rect 4375 31580 4439 31584
rect 4375 31524 4379 31580
rect 4379 31524 4435 31580
rect 4435 31524 4439 31580
rect 4375 31520 4439 31524
rect 4455 31580 4519 31584
rect 4455 31524 4459 31580
rect 4459 31524 4515 31580
rect 4515 31524 4519 31580
rect 4455 31520 4519 31524
rect 7479 31580 7543 31584
rect 7479 31524 7483 31580
rect 7483 31524 7539 31580
rect 7539 31524 7543 31580
rect 7479 31520 7543 31524
rect 7559 31580 7623 31584
rect 7559 31524 7563 31580
rect 7563 31524 7619 31580
rect 7619 31524 7623 31580
rect 7559 31520 7623 31524
rect 7639 31580 7703 31584
rect 7639 31524 7643 31580
rect 7643 31524 7699 31580
rect 7699 31524 7703 31580
rect 7639 31520 7703 31524
rect 7719 31580 7783 31584
rect 7719 31524 7723 31580
rect 7723 31524 7779 31580
rect 7779 31524 7783 31580
rect 7719 31520 7783 31524
rect 2584 31036 2648 31040
rect 2584 30980 2588 31036
rect 2588 30980 2644 31036
rect 2644 30980 2648 31036
rect 2584 30976 2648 30980
rect 2664 31036 2728 31040
rect 2664 30980 2668 31036
rect 2668 30980 2724 31036
rect 2724 30980 2728 31036
rect 2664 30976 2728 30980
rect 2744 31036 2808 31040
rect 2744 30980 2748 31036
rect 2748 30980 2804 31036
rect 2804 30980 2808 31036
rect 2744 30976 2808 30980
rect 2824 31036 2888 31040
rect 2824 30980 2828 31036
rect 2828 30980 2884 31036
rect 2884 30980 2888 31036
rect 2824 30976 2888 30980
rect 5847 31036 5911 31040
rect 5847 30980 5851 31036
rect 5851 30980 5907 31036
rect 5907 30980 5911 31036
rect 5847 30976 5911 30980
rect 5927 31036 5991 31040
rect 5927 30980 5931 31036
rect 5931 30980 5987 31036
rect 5987 30980 5991 31036
rect 5927 30976 5991 30980
rect 6007 31036 6071 31040
rect 6007 30980 6011 31036
rect 6011 30980 6067 31036
rect 6067 30980 6071 31036
rect 6007 30976 6071 30980
rect 6087 31036 6151 31040
rect 6087 30980 6091 31036
rect 6091 30980 6147 31036
rect 6147 30980 6151 31036
rect 6087 30976 6151 30980
rect 9111 31036 9175 31040
rect 9111 30980 9115 31036
rect 9115 30980 9171 31036
rect 9171 30980 9175 31036
rect 9111 30976 9175 30980
rect 9191 31036 9255 31040
rect 9191 30980 9195 31036
rect 9195 30980 9251 31036
rect 9251 30980 9255 31036
rect 9191 30976 9255 30980
rect 9271 31036 9335 31040
rect 9271 30980 9275 31036
rect 9275 30980 9331 31036
rect 9331 30980 9335 31036
rect 9271 30976 9335 30980
rect 9351 31036 9415 31040
rect 9351 30980 9355 31036
rect 9355 30980 9411 31036
rect 9411 30980 9415 31036
rect 9351 30976 9415 30980
rect 4215 30492 4279 30496
rect 4215 30436 4219 30492
rect 4219 30436 4275 30492
rect 4275 30436 4279 30492
rect 4215 30432 4279 30436
rect 4295 30492 4359 30496
rect 4295 30436 4299 30492
rect 4299 30436 4355 30492
rect 4355 30436 4359 30492
rect 4295 30432 4359 30436
rect 4375 30492 4439 30496
rect 4375 30436 4379 30492
rect 4379 30436 4435 30492
rect 4435 30436 4439 30492
rect 4375 30432 4439 30436
rect 4455 30492 4519 30496
rect 4455 30436 4459 30492
rect 4459 30436 4515 30492
rect 4515 30436 4519 30492
rect 4455 30432 4519 30436
rect 7479 30492 7543 30496
rect 7479 30436 7483 30492
rect 7483 30436 7539 30492
rect 7539 30436 7543 30492
rect 7479 30432 7543 30436
rect 7559 30492 7623 30496
rect 7559 30436 7563 30492
rect 7563 30436 7619 30492
rect 7619 30436 7623 30492
rect 7559 30432 7623 30436
rect 7639 30492 7703 30496
rect 7639 30436 7643 30492
rect 7643 30436 7699 30492
rect 7699 30436 7703 30492
rect 7639 30432 7703 30436
rect 7719 30492 7783 30496
rect 7719 30436 7723 30492
rect 7723 30436 7779 30492
rect 7779 30436 7783 30492
rect 7719 30432 7783 30436
rect 2584 29948 2648 29952
rect 2584 29892 2588 29948
rect 2588 29892 2644 29948
rect 2644 29892 2648 29948
rect 2584 29888 2648 29892
rect 2664 29948 2728 29952
rect 2664 29892 2668 29948
rect 2668 29892 2724 29948
rect 2724 29892 2728 29948
rect 2664 29888 2728 29892
rect 2744 29948 2808 29952
rect 2744 29892 2748 29948
rect 2748 29892 2804 29948
rect 2804 29892 2808 29948
rect 2744 29888 2808 29892
rect 2824 29948 2888 29952
rect 2824 29892 2828 29948
rect 2828 29892 2884 29948
rect 2884 29892 2888 29948
rect 2824 29888 2888 29892
rect 5847 29948 5911 29952
rect 5847 29892 5851 29948
rect 5851 29892 5907 29948
rect 5907 29892 5911 29948
rect 5847 29888 5911 29892
rect 5927 29948 5991 29952
rect 5927 29892 5931 29948
rect 5931 29892 5987 29948
rect 5987 29892 5991 29948
rect 5927 29888 5991 29892
rect 6007 29948 6071 29952
rect 6007 29892 6011 29948
rect 6011 29892 6067 29948
rect 6067 29892 6071 29948
rect 6007 29888 6071 29892
rect 6087 29948 6151 29952
rect 6087 29892 6091 29948
rect 6091 29892 6147 29948
rect 6147 29892 6151 29948
rect 6087 29888 6151 29892
rect 9111 29948 9175 29952
rect 9111 29892 9115 29948
rect 9115 29892 9171 29948
rect 9171 29892 9175 29948
rect 9111 29888 9175 29892
rect 9191 29948 9255 29952
rect 9191 29892 9195 29948
rect 9195 29892 9251 29948
rect 9251 29892 9255 29948
rect 9191 29888 9255 29892
rect 9271 29948 9335 29952
rect 9271 29892 9275 29948
rect 9275 29892 9331 29948
rect 9331 29892 9335 29948
rect 9271 29888 9335 29892
rect 9351 29948 9415 29952
rect 9351 29892 9355 29948
rect 9355 29892 9411 29948
rect 9411 29892 9415 29948
rect 9351 29888 9415 29892
rect 4215 29404 4279 29408
rect 4215 29348 4219 29404
rect 4219 29348 4275 29404
rect 4275 29348 4279 29404
rect 4215 29344 4279 29348
rect 4295 29404 4359 29408
rect 4295 29348 4299 29404
rect 4299 29348 4355 29404
rect 4355 29348 4359 29404
rect 4295 29344 4359 29348
rect 4375 29404 4439 29408
rect 4375 29348 4379 29404
rect 4379 29348 4435 29404
rect 4435 29348 4439 29404
rect 4375 29344 4439 29348
rect 4455 29404 4519 29408
rect 4455 29348 4459 29404
rect 4459 29348 4515 29404
rect 4515 29348 4519 29404
rect 4455 29344 4519 29348
rect 7479 29404 7543 29408
rect 7479 29348 7483 29404
rect 7483 29348 7539 29404
rect 7539 29348 7543 29404
rect 7479 29344 7543 29348
rect 7559 29404 7623 29408
rect 7559 29348 7563 29404
rect 7563 29348 7619 29404
rect 7619 29348 7623 29404
rect 7559 29344 7623 29348
rect 7639 29404 7703 29408
rect 7639 29348 7643 29404
rect 7643 29348 7699 29404
rect 7699 29348 7703 29404
rect 7639 29344 7703 29348
rect 7719 29404 7783 29408
rect 7719 29348 7723 29404
rect 7723 29348 7779 29404
rect 7779 29348 7783 29404
rect 7719 29344 7783 29348
rect 2584 28860 2648 28864
rect 2584 28804 2588 28860
rect 2588 28804 2644 28860
rect 2644 28804 2648 28860
rect 2584 28800 2648 28804
rect 2664 28860 2728 28864
rect 2664 28804 2668 28860
rect 2668 28804 2724 28860
rect 2724 28804 2728 28860
rect 2664 28800 2728 28804
rect 2744 28860 2808 28864
rect 2744 28804 2748 28860
rect 2748 28804 2804 28860
rect 2804 28804 2808 28860
rect 2744 28800 2808 28804
rect 2824 28860 2888 28864
rect 2824 28804 2828 28860
rect 2828 28804 2884 28860
rect 2884 28804 2888 28860
rect 2824 28800 2888 28804
rect 5847 28860 5911 28864
rect 5847 28804 5851 28860
rect 5851 28804 5907 28860
rect 5907 28804 5911 28860
rect 5847 28800 5911 28804
rect 5927 28860 5991 28864
rect 5927 28804 5931 28860
rect 5931 28804 5987 28860
rect 5987 28804 5991 28860
rect 5927 28800 5991 28804
rect 6007 28860 6071 28864
rect 6007 28804 6011 28860
rect 6011 28804 6067 28860
rect 6067 28804 6071 28860
rect 6007 28800 6071 28804
rect 6087 28860 6151 28864
rect 6087 28804 6091 28860
rect 6091 28804 6147 28860
rect 6147 28804 6151 28860
rect 6087 28800 6151 28804
rect 9111 28860 9175 28864
rect 9111 28804 9115 28860
rect 9115 28804 9171 28860
rect 9171 28804 9175 28860
rect 9111 28800 9175 28804
rect 9191 28860 9255 28864
rect 9191 28804 9195 28860
rect 9195 28804 9251 28860
rect 9251 28804 9255 28860
rect 9191 28800 9255 28804
rect 9271 28860 9335 28864
rect 9271 28804 9275 28860
rect 9275 28804 9331 28860
rect 9331 28804 9335 28860
rect 9271 28800 9335 28804
rect 9351 28860 9415 28864
rect 9351 28804 9355 28860
rect 9355 28804 9411 28860
rect 9411 28804 9415 28860
rect 9351 28800 9415 28804
rect 4215 28316 4279 28320
rect 4215 28260 4219 28316
rect 4219 28260 4275 28316
rect 4275 28260 4279 28316
rect 4215 28256 4279 28260
rect 4295 28316 4359 28320
rect 4295 28260 4299 28316
rect 4299 28260 4355 28316
rect 4355 28260 4359 28316
rect 4295 28256 4359 28260
rect 4375 28316 4439 28320
rect 4375 28260 4379 28316
rect 4379 28260 4435 28316
rect 4435 28260 4439 28316
rect 4375 28256 4439 28260
rect 4455 28316 4519 28320
rect 4455 28260 4459 28316
rect 4459 28260 4515 28316
rect 4515 28260 4519 28316
rect 4455 28256 4519 28260
rect 7479 28316 7543 28320
rect 7479 28260 7483 28316
rect 7483 28260 7539 28316
rect 7539 28260 7543 28316
rect 7479 28256 7543 28260
rect 7559 28316 7623 28320
rect 7559 28260 7563 28316
rect 7563 28260 7619 28316
rect 7619 28260 7623 28316
rect 7559 28256 7623 28260
rect 7639 28316 7703 28320
rect 7639 28260 7643 28316
rect 7643 28260 7699 28316
rect 7699 28260 7703 28316
rect 7639 28256 7703 28260
rect 7719 28316 7783 28320
rect 7719 28260 7723 28316
rect 7723 28260 7779 28316
rect 7779 28260 7783 28316
rect 7719 28256 7783 28260
rect 2584 27772 2648 27776
rect 2584 27716 2588 27772
rect 2588 27716 2644 27772
rect 2644 27716 2648 27772
rect 2584 27712 2648 27716
rect 2664 27772 2728 27776
rect 2664 27716 2668 27772
rect 2668 27716 2724 27772
rect 2724 27716 2728 27772
rect 2664 27712 2728 27716
rect 2744 27772 2808 27776
rect 2744 27716 2748 27772
rect 2748 27716 2804 27772
rect 2804 27716 2808 27772
rect 2744 27712 2808 27716
rect 2824 27772 2888 27776
rect 2824 27716 2828 27772
rect 2828 27716 2884 27772
rect 2884 27716 2888 27772
rect 2824 27712 2888 27716
rect 5847 27772 5911 27776
rect 5847 27716 5851 27772
rect 5851 27716 5907 27772
rect 5907 27716 5911 27772
rect 5847 27712 5911 27716
rect 5927 27772 5991 27776
rect 5927 27716 5931 27772
rect 5931 27716 5987 27772
rect 5987 27716 5991 27772
rect 5927 27712 5991 27716
rect 6007 27772 6071 27776
rect 6007 27716 6011 27772
rect 6011 27716 6067 27772
rect 6067 27716 6071 27772
rect 6007 27712 6071 27716
rect 6087 27772 6151 27776
rect 6087 27716 6091 27772
rect 6091 27716 6147 27772
rect 6147 27716 6151 27772
rect 6087 27712 6151 27716
rect 9111 27772 9175 27776
rect 9111 27716 9115 27772
rect 9115 27716 9171 27772
rect 9171 27716 9175 27772
rect 9111 27712 9175 27716
rect 9191 27772 9255 27776
rect 9191 27716 9195 27772
rect 9195 27716 9251 27772
rect 9251 27716 9255 27772
rect 9191 27712 9255 27716
rect 9271 27772 9335 27776
rect 9271 27716 9275 27772
rect 9275 27716 9331 27772
rect 9331 27716 9335 27772
rect 9271 27712 9335 27716
rect 9351 27772 9415 27776
rect 9351 27716 9355 27772
rect 9355 27716 9411 27772
rect 9411 27716 9415 27772
rect 9351 27712 9415 27716
rect 4215 27228 4279 27232
rect 4215 27172 4219 27228
rect 4219 27172 4275 27228
rect 4275 27172 4279 27228
rect 4215 27168 4279 27172
rect 4295 27228 4359 27232
rect 4295 27172 4299 27228
rect 4299 27172 4355 27228
rect 4355 27172 4359 27228
rect 4295 27168 4359 27172
rect 4375 27228 4439 27232
rect 4375 27172 4379 27228
rect 4379 27172 4435 27228
rect 4435 27172 4439 27228
rect 4375 27168 4439 27172
rect 4455 27228 4519 27232
rect 4455 27172 4459 27228
rect 4459 27172 4515 27228
rect 4515 27172 4519 27228
rect 4455 27168 4519 27172
rect 7479 27228 7543 27232
rect 7479 27172 7483 27228
rect 7483 27172 7539 27228
rect 7539 27172 7543 27228
rect 7479 27168 7543 27172
rect 7559 27228 7623 27232
rect 7559 27172 7563 27228
rect 7563 27172 7619 27228
rect 7619 27172 7623 27228
rect 7559 27168 7623 27172
rect 7639 27228 7703 27232
rect 7639 27172 7643 27228
rect 7643 27172 7699 27228
rect 7699 27172 7703 27228
rect 7639 27168 7703 27172
rect 7719 27228 7783 27232
rect 7719 27172 7723 27228
rect 7723 27172 7779 27228
rect 7779 27172 7783 27228
rect 7719 27168 7783 27172
rect 2584 26684 2648 26688
rect 2584 26628 2588 26684
rect 2588 26628 2644 26684
rect 2644 26628 2648 26684
rect 2584 26624 2648 26628
rect 2664 26684 2728 26688
rect 2664 26628 2668 26684
rect 2668 26628 2724 26684
rect 2724 26628 2728 26684
rect 2664 26624 2728 26628
rect 2744 26684 2808 26688
rect 2744 26628 2748 26684
rect 2748 26628 2804 26684
rect 2804 26628 2808 26684
rect 2744 26624 2808 26628
rect 2824 26684 2888 26688
rect 2824 26628 2828 26684
rect 2828 26628 2884 26684
rect 2884 26628 2888 26684
rect 2824 26624 2888 26628
rect 5847 26684 5911 26688
rect 5847 26628 5851 26684
rect 5851 26628 5907 26684
rect 5907 26628 5911 26684
rect 5847 26624 5911 26628
rect 5927 26684 5991 26688
rect 5927 26628 5931 26684
rect 5931 26628 5987 26684
rect 5987 26628 5991 26684
rect 5927 26624 5991 26628
rect 6007 26684 6071 26688
rect 6007 26628 6011 26684
rect 6011 26628 6067 26684
rect 6067 26628 6071 26684
rect 6007 26624 6071 26628
rect 6087 26684 6151 26688
rect 6087 26628 6091 26684
rect 6091 26628 6147 26684
rect 6147 26628 6151 26684
rect 6087 26624 6151 26628
rect 9111 26684 9175 26688
rect 9111 26628 9115 26684
rect 9115 26628 9171 26684
rect 9171 26628 9175 26684
rect 9111 26624 9175 26628
rect 9191 26684 9255 26688
rect 9191 26628 9195 26684
rect 9195 26628 9251 26684
rect 9251 26628 9255 26684
rect 9191 26624 9255 26628
rect 9271 26684 9335 26688
rect 9271 26628 9275 26684
rect 9275 26628 9331 26684
rect 9331 26628 9335 26684
rect 9271 26624 9335 26628
rect 9351 26684 9415 26688
rect 9351 26628 9355 26684
rect 9355 26628 9411 26684
rect 9411 26628 9415 26684
rect 9351 26624 9415 26628
rect 4215 26140 4279 26144
rect 4215 26084 4219 26140
rect 4219 26084 4275 26140
rect 4275 26084 4279 26140
rect 4215 26080 4279 26084
rect 4295 26140 4359 26144
rect 4295 26084 4299 26140
rect 4299 26084 4355 26140
rect 4355 26084 4359 26140
rect 4295 26080 4359 26084
rect 4375 26140 4439 26144
rect 4375 26084 4379 26140
rect 4379 26084 4435 26140
rect 4435 26084 4439 26140
rect 4375 26080 4439 26084
rect 4455 26140 4519 26144
rect 4455 26084 4459 26140
rect 4459 26084 4515 26140
rect 4515 26084 4519 26140
rect 4455 26080 4519 26084
rect 7479 26140 7543 26144
rect 7479 26084 7483 26140
rect 7483 26084 7539 26140
rect 7539 26084 7543 26140
rect 7479 26080 7543 26084
rect 7559 26140 7623 26144
rect 7559 26084 7563 26140
rect 7563 26084 7619 26140
rect 7619 26084 7623 26140
rect 7559 26080 7623 26084
rect 7639 26140 7703 26144
rect 7639 26084 7643 26140
rect 7643 26084 7699 26140
rect 7699 26084 7703 26140
rect 7639 26080 7703 26084
rect 7719 26140 7783 26144
rect 7719 26084 7723 26140
rect 7723 26084 7779 26140
rect 7779 26084 7783 26140
rect 7719 26080 7783 26084
rect 2584 25596 2648 25600
rect 2584 25540 2588 25596
rect 2588 25540 2644 25596
rect 2644 25540 2648 25596
rect 2584 25536 2648 25540
rect 2664 25596 2728 25600
rect 2664 25540 2668 25596
rect 2668 25540 2724 25596
rect 2724 25540 2728 25596
rect 2664 25536 2728 25540
rect 2744 25596 2808 25600
rect 2744 25540 2748 25596
rect 2748 25540 2804 25596
rect 2804 25540 2808 25596
rect 2744 25536 2808 25540
rect 2824 25596 2888 25600
rect 2824 25540 2828 25596
rect 2828 25540 2884 25596
rect 2884 25540 2888 25596
rect 2824 25536 2888 25540
rect 5847 25596 5911 25600
rect 5847 25540 5851 25596
rect 5851 25540 5907 25596
rect 5907 25540 5911 25596
rect 5847 25536 5911 25540
rect 5927 25596 5991 25600
rect 5927 25540 5931 25596
rect 5931 25540 5987 25596
rect 5987 25540 5991 25596
rect 5927 25536 5991 25540
rect 6007 25596 6071 25600
rect 6007 25540 6011 25596
rect 6011 25540 6067 25596
rect 6067 25540 6071 25596
rect 6007 25536 6071 25540
rect 6087 25596 6151 25600
rect 6087 25540 6091 25596
rect 6091 25540 6147 25596
rect 6147 25540 6151 25596
rect 6087 25536 6151 25540
rect 9111 25596 9175 25600
rect 9111 25540 9115 25596
rect 9115 25540 9171 25596
rect 9171 25540 9175 25596
rect 9111 25536 9175 25540
rect 9191 25596 9255 25600
rect 9191 25540 9195 25596
rect 9195 25540 9251 25596
rect 9251 25540 9255 25596
rect 9191 25536 9255 25540
rect 9271 25596 9335 25600
rect 9271 25540 9275 25596
rect 9275 25540 9331 25596
rect 9331 25540 9335 25596
rect 9271 25536 9335 25540
rect 9351 25596 9415 25600
rect 9351 25540 9355 25596
rect 9355 25540 9411 25596
rect 9411 25540 9415 25596
rect 9351 25536 9415 25540
rect 4215 25052 4279 25056
rect 4215 24996 4219 25052
rect 4219 24996 4275 25052
rect 4275 24996 4279 25052
rect 4215 24992 4279 24996
rect 4295 25052 4359 25056
rect 4295 24996 4299 25052
rect 4299 24996 4355 25052
rect 4355 24996 4359 25052
rect 4295 24992 4359 24996
rect 4375 25052 4439 25056
rect 4375 24996 4379 25052
rect 4379 24996 4435 25052
rect 4435 24996 4439 25052
rect 4375 24992 4439 24996
rect 4455 25052 4519 25056
rect 4455 24996 4459 25052
rect 4459 24996 4515 25052
rect 4515 24996 4519 25052
rect 4455 24992 4519 24996
rect 7479 25052 7543 25056
rect 7479 24996 7483 25052
rect 7483 24996 7539 25052
rect 7539 24996 7543 25052
rect 7479 24992 7543 24996
rect 7559 25052 7623 25056
rect 7559 24996 7563 25052
rect 7563 24996 7619 25052
rect 7619 24996 7623 25052
rect 7559 24992 7623 24996
rect 7639 25052 7703 25056
rect 7639 24996 7643 25052
rect 7643 24996 7699 25052
rect 7699 24996 7703 25052
rect 7639 24992 7703 24996
rect 7719 25052 7783 25056
rect 7719 24996 7723 25052
rect 7723 24996 7779 25052
rect 7779 24996 7783 25052
rect 7719 24992 7783 24996
rect 2584 24508 2648 24512
rect 2584 24452 2588 24508
rect 2588 24452 2644 24508
rect 2644 24452 2648 24508
rect 2584 24448 2648 24452
rect 2664 24508 2728 24512
rect 2664 24452 2668 24508
rect 2668 24452 2724 24508
rect 2724 24452 2728 24508
rect 2664 24448 2728 24452
rect 2744 24508 2808 24512
rect 2744 24452 2748 24508
rect 2748 24452 2804 24508
rect 2804 24452 2808 24508
rect 2744 24448 2808 24452
rect 2824 24508 2888 24512
rect 2824 24452 2828 24508
rect 2828 24452 2884 24508
rect 2884 24452 2888 24508
rect 2824 24448 2888 24452
rect 5847 24508 5911 24512
rect 5847 24452 5851 24508
rect 5851 24452 5907 24508
rect 5907 24452 5911 24508
rect 5847 24448 5911 24452
rect 5927 24508 5991 24512
rect 5927 24452 5931 24508
rect 5931 24452 5987 24508
rect 5987 24452 5991 24508
rect 5927 24448 5991 24452
rect 6007 24508 6071 24512
rect 6007 24452 6011 24508
rect 6011 24452 6067 24508
rect 6067 24452 6071 24508
rect 6007 24448 6071 24452
rect 6087 24508 6151 24512
rect 6087 24452 6091 24508
rect 6091 24452 6147 24508
rect 6147 24452 6151 24508
rect 6087 24448 6151 24452
rect 9111 24508 9175 24512
rect 9111 24452 9115 24508
rect 9115 24452 9171 24508
rect 9171 24452 9175 24508
rect 9111 24448 9175 24452
rect 9191 24508 9255 24512
rect 9191 24452 9195 24508
rect 9195 24452 9251 24508
rect 9251 24452 9255 24508
rect 9191 24448 9255 24452
rect 9271 24508 9335 24512
rect 9271 24452 9275 24508
rect 9275 24452 9331 24508
rect 9331 24452 9335 24508
rect 9271 24448 9335 24452
rect 9351 24508 9415 24512
rect 9351 24452 9355 24508
rect 9355 24452 9411 24508
rect 9411 24452 9415 24508
rect 9351 24448 9415 24452
rect 4215 23964 4279 23968
rect 4215 23908 4219 23964
rect 4219 23908 4275 23964
rect 4275 23908 4279 23964
rect 4215 23904 4279 23908
rect 4295 23964 4359 23968
rect 4295 23908 4299 23964
rect 4299 23908 4355 23964
rect 4355 23908 4359 23964
rect 4295 23904 4359 23908
rect 4375 23964 4439 23968
rect 4375 23908 4379 23964
rect 4379 23908 4435 23964
rect 4435 23908 4439 23964
rect 4375 23904 4439 23908
rect 4455 23964 4519 23968
rect 4455 23908 4459 23964
rect 4459 23908 4515 23964
rect 4515 23908 4519 23964
rect 4455 23904 4519 23908
rect 7479 23964 7543 23968
rect 7479 23908 7483 23964
rect 7483 23908 7539 23964
rect 7539 23908 7543 23964
rect 7479 23904 7543 23908
rect 7559 23964 7623 23968
rect 7559 23908 7563 23964
rect 7563 23908 7619 23964
rect 7619 23908 7623 23964
rect 7559 23904 7623 23908
rect 7639 23964 7703 23968
rect 7639 23908 7643 23964
rect 7643 23908 7699 23964
rect 7699 23908 7703 23964
rect 7639 23904 7703 23908
rect 7719 23964 7783 23968
rect 7719 23908 7723 23964
rect 7723 23908 7779 23964
rect 7779 23908 7783 23964
rect 7719 23904 7783 23908
rect 2584 23420 2648 23424
rect 2584 23364 2588 23420
rect 2588 23364 2644 23420
rect 2644 23364 2648 23420
rect 2584 23360 2648 23364
rect 2664 23420 2728 23424
rect 2664 23364 2668 23420
rect 2668 23364 2724 23420
rect 2724 23364 2728 23420
rect 2664 23360 2728 23364
rect 2744 23420 2808 23424
rect 2744 23364 2748 23420
rect 2748 23364 2804 23420
rect 2804 23364 2808 23420
rect 2744 23360 2808 23364
rect 2824 23420 2888 23424
rect 2824 23364 2828 23420
rect 2828 23364 2884 23420
rect 2884 23364 2888 23420
rect 2824 23360 2888 23364
rect 5847 23420 5911 23424
rect 5847 23364 5851 23420
rect 5851 23364 5907 23420
rect 5907 23364 5911 23420
rect 5847 23360 5911 23364
rect 5927 23420 5991 23424
rect 5927 23364 5931 23420
rect 5931 23364 5987 23420
rect 5987 23364 5991 23420
rect 5927 23360 5991 23364
rect 6007 23420 6071 23424
rect 6007 23364 6011 23420
rect 6011 23364 6067 23420
rect 6067 23364 6071 23420
rect 6007 23360 6071 23364
rect 6087 23420 6151 23424
rect 6087 23364 6091 23420
rect 6091 23364 6147 23420
rect 6147 23364 6151 23420
rect 6087 23360 6151 23364
rect 9111 23420 9175 23424
rect 9111 23364 9115 23420
rect 9115 23364 9171 23420
rect 9171 23364 9175 23420
rect 9111 23360 9175 23364
rect 9191 23420 9255 23424
rect 9191 23364 9195 23420
rect 9195 23364 9251 23420
rect 9251 23364 9255 23420
rect 9191 23360 9255 23364
rect 9271 23420 9335 23424
rect 9271 23364 9275 23420
rect 9275 23364 9331 23420
rect 9331 23364 9335 23420
rect 9271 23360 9335 23364
rect 9351 23420 9415 23424
rect 9351 23364 9355 23420
rect 9355 23364 9411 23420
rect 9411 23364 9415 23420
rect 9351 23360 9415 23364
rect 4215 22876 4279 22880
rect 4215 22820 4219 22876
rect 4219 22820 4275 22876
rect 4275 22820 4279 22876
rect 4215 22816 4279 22820
rect 4295 22876 4359 22880
rect 4295 22820 4299 22876
rect 4299 22820 4355 22876
rect 4355 22820 4359 22876
rect 4295 22816 4359 22820
rect 4375 22876 4439 22880
rect 4375 22820 4379 22876
rect 4379 22820 4435 22876
rect 4435 22820 4439 22876
rect 4375 22816 4439 22820
rect 4455 22876 4519 22880
rect 4455 22820 4459 22876
rect 4459 22820 4515 22876
rect 4515 22820 4519 22876
rect 4455 22816 4519 22820
rect 7479 22876 7543 22880
rect 7479 22820 7483 22876
rect 7483 22820 7539 22876
rect 7539 22820 7543 22876
rect 7479 22816 7543 22820
rect 7559 22876 7623 22880
rect 7559 22820 7563 22876
rect 7563 22820 7619 22876
rect 7619 22820 7623 22876
rect 7559 22816 7623 22820
rect 7639 22876 7703 22880
rect 7639 22820 7643 22876
rect 7643 22820 7699 22876
rect 7699 22820 7703 22876
rect 7639 22816 7703 22820
rect 7719 22876 7783 22880
rect 7719 22820 7723 22876
rect 7723 22820 7779 22876
rect 7779 22820 7783 22876
rect 7719 22816 7783 22820
rect 2584 22332 2648 22336
rect 2584 22276 2588 22332
rect 2588 22276 2644 22332
rect 2644 22276 2648 22332
rect 2584 22272 2648 22276
rect 2664 22332 2728 22336
rect 2664 22276 2668 22332
rect 2668 22276 2724 22332
rect 2724 22276 2728 22332
rect 2664 22272 2728 22276
rect 2744 22332 2808 22336
rect 2744 22276 2748 22332
rect 2748 22276 2804 22332
rect 2804 22276 2808 22332
rect 2744 22272 2808 22276
rect 2824 22332 2888 22336
rect 2824 22276 2828 22332
rect 2828 22276 2884 22332
rect 2884 22276 2888 22332
rect 2824 22272 2888 22276
rect 5847 22332 5911 22336
rect 5847 22276 5851 22332
rect 5851 22276 5907 22332
rect 5907 22276 5911 22332
rect 5847 22272 5911 22276
rect 5927 22332 5991 22336
rect 5927 22276 5931 22332
rect 5931 22276 5987 22332
rect 5987 22276 5991 22332
rect 5927 22272 5991 22276
rect 6007 22332 6071 22336
rect 6007 22276 6011 22332
rect 6011 22276 6067 22332
rect 6067 22276 6071 22332
rect 6007 22272 6071 22276
rect 6087 22332 6151 22336
rect 6087 22276 6091 22332
rect 6091 22276 6147 22332
rect 6147 22276 6151 22332
rect 6087 22272 6151 22276
rect 9111 22332 9175 22336
rect 9111 22276 9115 22332
rect 9115 22276 9171 22332
rect 9171 22276 9175 22332
rect 9111 22272 9175 22276
rect 9191 22332 9255 22336
rect 9191 22276 9195 22332
rect 9195 22276 9251 22332
rect 9251 22276 9255 22332
rect 9191 22272 9255 22276
rect 9271 22332 9335 22336
rect 9271 22276 9275 22332
rect 9275 22276 9331 22332
rect 9331 22276 9335 22332
rect 9271 22272 9335 22276
rect 9351 22332 9415 22336
rect 9351 22276 9355 22332
rect 9355 22276 9411 22332
rect 9411 22276 9415 22332
rect 9351 22272 9415 22276
rect 4215 21788 4279 21792
rect 4215 21732 4219 21788
rect 4219 21732 4275 21788
rect 4275 21732 4279 21788
rect 4215 21728 4279 21732
rect 4295 21788 4359 21792
rect 4295 21732 4299 21788
rect 4299 21732 4355 21788
rect 4355 21732 4359 21788
rect 4295 21728 4359 21732
rect 4375 21788 4439 21792
rect 4375 21732 4379 21788
rect 4379 21732 4435 21788
rect 4435 21732 4439 21788
rect 4375 21728 4439 21732
rect 4455 21788 4519 21792
rect 4455 21732 4459 21788
rect 4459 21732 4515 21788
rect 4515 21732 4519 21788
rect 4455 21728 4519 21732
rect 7479 21788 7543 21792
rect 7479 21732 7483 21788
rect 7483 21732 7539 21788
rect 7539 21732 7543 21788
rect 7479 21728 7543 21732
rect 7559 21788 7623 21792
rect 7559 21732 7563 21788
rect 7563 21732 7619 21788
rect 7619 21732 7623 21788
rect 7559 21728 7623 21732
rect 7639 21788 7703 21792
rect 7639 21732 7643 21788
rect 7643 21732 7699 21788
rect 7699 21732 7703 21788
rect 7639 21728 7703 21732
rect 7719 21788 7783 21792
rect 7719 21732 7723 21788
rect 7723 21732 7779 21788
rect 7779 21732 7783 21788
rect 7719 21728 7783 21732
rect 2584 21244 2648 21248
rect 2584 21188 2588 21244
rect 2588 21188 2644 21244
rect 2644 21188 2648 21244
rect 2584 21184 2648 21188
rect 2664 21244 2728 21248
rect 2664 21188 2668 21244
rect 2668 21188 2724 21244
rect 2724 21188 2728 21244
rect 2664 21184 2728 21188
rect 2744 21244 2808 21248
rect 2744 21188 2748 21244
rect 2748 21188 2804 21244
rect 2804 21188 2808 21244
rect 2744 21184 2808 21188
rect 2824 21244 2888 21248
rect 2824 21188 2828 21244
rect 2828 21188 2884 21244
rect 2884 21188 2888 21244
rect 2824 21184 2888 21188
rect 5847 21244 5911 21248
rect 5847 21188 5851 21244
rect 5851 21188 5907 21244
rect 5907 21188 5911 21244
rect 5847 21184 5911 21188
rect 5927 21244 5991 21248
rect 5927 21188 5931 21244
rect 5931 21188 5987 21244
rect 5987 21188 5991 21244
rect 5927 21184 5991 21188
rect 6007 21244 6071 21248
rect 6007 21188 6011 21244
rect 6011 21188 6067 21244
rect 6067 21188 6071 21244
rect 6007 21184 6071 21188
rect 6087 21244 6151 21248
rect 6087 21188 6091 21244
rect 6091 21188 6147 21244
rect 6147 21188 6151 21244
rect 6087 21184 6151 21188
rect 9111 21244 9175 21248
rect 9111 21188 9115 21244
rect 9115 21188 9171 21244
rect 9171 21188 9175 21244
rect 9111 21184 9175 21188
rect 9191 21244 9255 21248
rect 9191 21188 9195 21244
rect 9195 21188 9251 21244
rect 9251 21188 9255 21244
rect 9191 21184 9255 21188
rect 9271 21244 9335 21248
rect 9271 21188 9275 21244
rect 9275 21188 9331 21244
rect 9331 21188 9335 21244
rect 9271 21184 9335 21188
rect 9351 21244 9415 21248
rect 9351 21188 9355 21244
rect 9355 21188 9411 21244
rect 9411 21188 9415 21244
rect 9351 21184 9415 21188
rect 4215 20700 4279 20704
rect 4215 20644 4219 20700
rect 4219 20644 4275 20700
rect 4275 20644 4279 20700
rect 4215 20640 4279 20644
rect 4295 20700 4359 20704
rect 4295 20644 4299 20700
rect 4299 20644 4355 20700
rect 4355 20644 4359 20700
rect 4295 20640 4359 20644
rect 4375 20700 4439 20704
rect 4375 20644 4379 20700
rect 4379 20644 4435 20700
rect 4435 20644 4439 20700
rect 4375 20640 4439 20644
rect 4455 20700 4519 20704
rect 4455 20644 4459 20700
rect 4459 20644 4515 20700
rect 4515 20644 4519 20700
rect 4455 20640 4519 20644
rect 7479 20700 7543 20704
rect 7479 20644 7483 20700
rect 7483 20644 7539 20700
rect 7539 20644 7543 20700
rect 7479 20640 7543 20644
rect 7559 20700 7623 20704
rect 7559 20644 7563 20700
rect 7563 20644 7619 20700
rect 7619 20644 7623 20700
rect 7559 20640 7623 20644
rect 7639 20700 7703 20704
rect 7639 20644 7643 20700
rect 7643 20644 7699 20700
rect 7699 20644 7703 20700
rect 7639 20640 7703 20644
rect 7719 20700 7783 20704
rect 7719 20644 7723 20700
rect 7723 20644 7779 20700
rect 7779 20644 7783 20700
rect 7719 20640 7783 20644
rect 2584 20156 2648 20160
rect 2584 20100 2588 20156
rect 2588 20100 2644 20156
rect 2644 20100 2648 20156
rect 2584 20096 2648 20100
rect 2664 20156 2728 20160
rect 2664 20100 2668 20156
rect 2668 20100 2724 20156
rect 2724 20100 2728 20156
rect 2664 20096 2728 20100
rect 2744 20156 2808 20160
rect 2744 20100 2748 20156
rect 2748 20100 2804 20156
rect 2804 20100 2808 20156
rect 2744 20096 2808 20100
rect 2824 20156 2888 20160
rect 2824 20100 2828 20156
rect 2828 20100 2884 20156
rect 2884 20100 2888 20156
rect 2824 20096 2888 20100
rect 5847 20156 5911 20160
rect 5847 20100 5851 20156
rect 5851 20100 5907 20156
rect 5907 20100 5911 20156
rect 5847 20096 5911 20100
rect 5927 20156 5991 20160
rect 5927 20100 5931 20156
rect 5931 20100 5987 20156
rect 5987 20100 5991 20156
rect 5927 20096 5991 20100
rect 6007 20156 6071 20160
rect 6007 20100 6011 20156
rect 6011 20100 6067 20156
rect 6067 20100 6071 20156
rect 6007 20096 6071 20100
rect 6087 20156 6151 20160
rect 6087 20100 6091 20156
rect 6091 20100 6147 20156
rect 6147 20100 6151 20156
rect 6087 20096 6151 20100
rect 9111 20156 9175 20160
rect 9111 20100 9115 20156
rect 9115 20100 9171 20156
rect 9171 20100 9175 20156
rect 9111 20096 9175 20100
rect 9191 20156 9255 20160
rect 9191 20100 9195 20156
rect 9195 20100 9251 20156
rect 9251 20100 9255 20156
rect 9191 20096 9255 20100
rect 9271 20156 9335 20160
rect 9271 20100 9275 20156
rect 9275 20100 9331 20156
rect 9331 20100 9335 20156
rect 9271 20096 9335 20100
rect 9351 20156 9415 20160
rect 9351 20100 9355 20156
rect 9355 20100 9411 20156
rect 9411 20100 9415 20156
rect 9351 20096 9415 20100
rect 4215 19612 4279 19616
rect 4215 19556 4219 19612
rect 4219 19556 4275 19612
rect 4275 19556 4279 19612
rect 4215 19552 4279 19556
rect 4295 19612 4359 19616
rect 4295 19556 4299 19612
rect 4299 19556 4355 19612
rect 4355 19556 4359 19612
rect 4295 19552 4359 19556
rect 4375 19612 4439 19616
rect 4375 19556 4379 19612
rect 4379 19556 4435 19612
rect 4435 19556 4439 19612
rect 4375 19552 4439 19556
rect 4455 19612 4519 19616
rect 4455 19556 4459 19612
rect 4459 19556 4515 19612
rect 4515 19556 4519 19612
rect 4455 19552 4519 19556
rect 7479 19612 7543 19616
rect 7479 19556 7483 19612
rect 7483 19556 7539 19612
rect 7539 19556 7543 19612
rect 7479 19552 7543 19556
rect 7559 19612 7623 19616
rect 7559 19556 7563 19612
rect 7563 19556 7619 19612
rect 7619 19556 7623 19612
rect 7559 19552 7623 19556
rect 7639 19612 7703 19616
rect 7639 19556 7643 19612
rect 7643 19556 7699 19612
rect 7699 19556 7703 19612
rect 7639 19552 7703 19556
rect 7719 19612 7783 19616
rect 7719 19556 7723 19612
rect 7723 19556 7779 19612
rect 7779 19556 7783 19612
rect 7719 19552 7783 19556
rect 2584 19068 2648 19072
rect 2584 19012 2588 19068
rect 2588 19012 2644 19068
rect 2644 19012 2648 19068
rect 2584 19008 2648 19012
rect 2664 19068 2728 19072
rect 2664 19012 2668 19068
rect 2668 19012 2724 19068
rect 2724 19012 2728 19068
rect 2664 19008 2728 19012
rect 2744 19068 2808 19072
rect 2744 19012 2748 19068
rect 2748 19012 2804 19068
rect 2804 19012 2808 19068
rect 2744 19008 2808 19012
rect 2824 19068 2888 19072
rect 2824 19012 2828 19068
rect 2828 19012 2884 19068
rect 2884 19012 2888 19068
rect 2824 19008 2888 19012
rect 5847 19068 5911 19072
rect 5847 19012 5851 19068
rect 5851 19012 5907 19068
rect 5907 19012 5911 19068
rect 5847 19008 5911 19012
rect 5927 19068 5991 19072
rect 5927 19012 5931 19068
rect 5931 19012 5987 19068
rect 5987 19012 5991 19068
rect 5927 19008 5991 19012
rect 6007 19068 6071 19072
rect 6007 19012 6011 19068
rect 6011 19012 6067 19068
rect 6067 19012 6071 19068
rect 6007 19008 6071 19012
rect 6087 19068 6151 19072
rect 6087 19012 6091 19068
rect 6091 19012 6147 19068
rect 6147 19012 6151 19068
rect 6087 19008 6151 19012
rect 9111 19068 9175 19072
rect 9111 19012 9115 19068
rect 9115 19012 9171 19068
rect 9171 19012 9175 19068
rect 9111 19008 9175 19012
rect 9191 19068 9255 19072
rect 9191 19012 9195 19068
rect 9195 19012 9251 19068
rect 9251 19012 9255 19068
rect 9191 19008 9255 19012
rect 9271 19068 9335 19072
rect 9271 19012 9275 19068
rect 9275 19012 9331 19068
rect 9331 19012 9335 19068
rect 9271 19008 9335 19012
rect 9351 19068 9415 19072
rect 9351 19012 9355 19068
rect 9355 19012 9411 19068
rect 9411 19012 9415 19068
rect 9351 19008 9415 19012
rect 4215 18524 4279 18528
rect 4215 18468 4219 18524
rect 4219 18468 4275 18524
rect 4275 18468 4279 18524
rect 4215 18464 4279 18468
rect 4295 18524 4359 18528
rect 4295 18468 4299 18524
rect 4299 18468 4355 18524
rect 4355 18468 4359 18524
rect 4295 18464 4359 18468
rect 4375 18524 4439 18528
rect 4375 18468 4379 18524
rect 4379 18468 4435 18524
rect 4435 18468 4439 18524
rect 4375 18464 4439 18468
rect 4455 18524 4519 18528
rect 4455 18468 4459 18524
rect 4459 18468 4515 18524
rect 4515 18468 4519 18524
rect 4455 18464 4519 18468
rect 7479 18524 7543 18528
rect 7479 18468 7483 18524
rect 7483 18468 7539 18524
rect 7539 18468 7543 18524
rect 7479 18464 7543 18468
rect 7559 18524 7623 18528
rect 7559 18468 7563 18524
rect 7563 18468 7619 18524
rect 7619 18468 7623 18524
rect 7559 18464 7623 18468
rect 7639 18524 7703 18528
rect 7639 18468 7643 18524
rect 7643 18468 7699 18524
rect 7699 18468 7703 18524
rect 7639 18464 7703 18468
rect 7719 18524 7783 18528
rect 7719 18468 7723 18524
rect 7723 18468 7779 18524
rect 7779 18468 7783 18524
rect 7719 18464 7783 18468
rect 2584 17980 2648 17984
rect 2584 17924 2588 17980
rect 2588 17924 2644 17980
rect 2644 17924 2648 17980
rect 2584 17920 2648 17924
rect 2664 17980 2728 17984
rect 2664 17924 2668 17980
rect 2668 17924 2724 17980
rect 2724 17924 2728 17980
rect 2664 17920 2728 17924
rect 2744 17980 2808 17984
rect 2744 17924 2748 17980
rect 2748 17924 2804 17980
rect 2804 17924 2808 17980
rect 2744 17920 2808 17924
rect 2824 17980 2888 17984
rect 2824 17924 2828 17980
rect 2828 17924 2884 17980
rect 2884 17924 2888 17980
rect 2824 17920 2888 17924
rect 5847 17980 5911 17984
rect 5847 17924 5851 17980
rect 5851 17924 5907 17980
rect 5907 17924 5911 17980
rect 5847 17920 5911 17924
rect 5927 17980 5991 17984
rect 5927 17924 5931 17980
rect 5931 17924 5987 17980
rect 5987 17924 5991 17980
rect 5927 17920 5991 17924
rect 6007 17980 6071 17984
rect 6007 17924 6011 17980
rect 6011 17924 6067 17980
rect 6067 17924 6071 17980
rect 6007 17920 6071 17924
rect 6087 17980 6151 17984
rect 6087 17924 6091 17980
rect 6091 17924 6147 17980
rect 6147 17924 6151 17980
rect 6087 17920 6151 17924
rect 9111 17980 9175 17984
rect 9111 17924 9115 17980
rect 9115 17924 9171 17980
rect 9171 17924 9175 17980
rect 9111 17920 9175 17924
rect 9191 17980 9255 17984
rect 9191 17924 9195 17980
rect 9195 17924 9251 17980
rect 9251 17924 9255 17980
rect 9191 17920 9255 17924
rect 9271 17980 9335 17984
rect 9271 17924 9275 17980
rect 9275 17924 9331 17980
rect 9331 17924 9335 17980
rect 9271 17920 9335 17924
rect 9351 17980 9415 17984
rect 9351 17924 9355 17980
rect 9355 17924 9411 17980
rect 9411 17924 9415 17980
rect 9351 17920 9415 17924
rect 4215 17436 4279 17440
rect 4215 17380 4219 17436
rect 4219 17380 4275 17436
rect 4275 17380 4279 17436
rect 4215 17376 4279 17380
rect 4295 17436 4359 17440
rect 4295 17380 4299 17436
rect 4299 17380 4355 17436
rect 4355 17380 4359 17436
rect 4295 17376 4359 17380
rect 4375 17436 4439 17440
rect 4375 17380 4379 17436
rect 4379 17380 4435 17436
rect 4435 17380 4439 17436
rect 4375 17376 4439 17380
rect 4455 17436 4519 17440
rect 4455 17380 4459 17436
rect 4459 17380 4515 17436
rect 4515 17380 4519 17436
rect 4455 17376 4519 17380
rect 7479 17436 7543 17440
rect 7479 17380 7483 17436
rect 7483 17380 7539 17436
rect 7539 17380 7543 17436
rect 7479 17376 7543 17380
rect 7559 17436 7623 17440
rect 7559 17380 7563 17436
rect 7563 17380 7619 17436
rect 7619 17380 7623 17436
rect 7559 17376 7623 17380
rect 7639 17436 7703 17440
rect 7639 17380 7643 17436
rect 7643 17380 7699 17436
rect 7699 17380 7703 17436
rect 7639 17376 7703 17380
rect 7719 17436 7783 17440
rect 7719 17380 7723 17436
rect 7723 17380 7779 17436
rect 7779 17380 7783 17436
rect 7719 17376 7783 17380
rect 2584 16892 2648 16896
rect 2584 16836 2588 16892
rect 2588 16836 2644 16892
rect 2644 16836 2648 16892
rect 2584 16832 2648 16836
rect 2664 16892 2728 16896
rect 2664 16836 2668 16892
rect 2668 16836 2724 16892
rect 2724 16836 2728 16892
rect 2664 16832 2728 16836
rect 2744 16892 2808 16896
rect 2744 16836 2748 16892
rect 2748 16836 2804 16892
rect 2804 16836 2808 16892
rect 2744 16832 2808 16836
rect 2824 16892 2888 16896
rect 2824 16836 2828 16892
rect 2828 16836 2884 16892
rect 2884 16836 2888 16892
rect 2824 16832 2888 16836
rect 5847 16892 5911 16896
rect 5847 16836 5851 16892
rect 5851 16836 5907 16892
rect 5907 16836 5911 16892
rect 5847 16832 5911 16836
rect 5927 16892 5991 16896
rect 5927 16836 5931 16892
rect 5931 16836 5987 16892
rect 5987 16836 5991 16892
rect 5927 16832 5991 16836
rect 6007 16892 6071 16896
rect 6007 16836 6011 16892
rect 6011 16836 6067 16892
rect 6067 16836 6071 16892
rect 6007 16832 6071 16836
rect 6087 16892 6151 16896
rect 6087 16836 6091 16892
rect 6091 16836 6147 16892
rect 6147 16836 6151 16892
rect 6087 16832 6151 16836
rect 9111 16892 9175 16896
rect 9111 16836 9115 16892
rect 9115 16836 9171 16892
rect 9171 16836 9175 16892
rect 9111 16832 9175 16836
rect 9191 16892 9255 16896
rect 9191 16836 9195 16892
rect 9195 16836 9251 16892
rect 9251 16836 9255 16892
rect 9191 16832 9255 16836
rect 9271 16892 9335 16896
rect 9271 16836 9275 16892
rect 9275 16836 9331 16892
rect 9331 16836 9335 16892
rect 9271 16832 9335 16836
rect 9351 16892 9415 16896
rect 9351 16836 9355 16892
rect 9355 16836 9411 16892
rect 9411 16836 9415 16892
rect 9351 16832 9415 16836
rect 4215 16348 4279 16352
rect 4215 16292 4219 16348
rect 4219 16292 4275 16348
rect 4275 16292 4279 16348
rect 4215 16288 4279 16292
rect 4295 16348 4359 16352
rect 4295 16292 4299 16348
rect 4299 16292 4355 16348
rect 4355 16292 4359 16348
rect 4295 16288 4359 16292
rect 4375 16348 4439 16352
rect 4375 16292 4379 16348
rect 4379 16292 4435 16348
rect 4435 16292 4439 16348
rect 4375 16288 4439 16292
rect 4455 16348 4519 16352
rect 4455 16292 4459 16348
rect 4459 16292 4515 16348
rect 4515 16292 4519 16348
rect 4455 16288 4519 16292
rect 7479 16348 7543 16352
rect 7479 16292 7483 16348
rect 7483 16292 7539 16348
rect 7539 16292 7543 16348
rect 7479 16288 7543 16292
rect 7559 16348 7623 16352
rect 7559 16292 7563 16348
rect 7563 16292 7619 16348
rect 7619 16292 7623 16348
rect 7559 16288 7623 16292
rect 7639 16348 7703 16352
rect 7639 16292 7643 16348
rect 7643 16292 7699 16348
rect 7699 16292 7703 16348
rect 7639 16288 7703 16292
rect 7719 16348 7783 16352
rect 7719 16292 7723 16348
rect 7723 16292 7779 16348
rect 7779 16292 7783 16348
rect 7719 16288 7783 16292
rect 2584 15804 2648 15808
rect 2584 15748 2588 15804
rect 2588 15748 2644 15804
rect 2644 15748 2648 15804
rect 2584 15744 2648 15748
rect 2664 15804 2728 15808
rect 2664 15748 2668 15804
rect 2668 15748 2724 15804
rect 2724 15748 2728 15804
rect 2664 15744 2728 15748
rect 2744 15804 2808 15808
rect 2744 15748 2748 15804
rect 2748 15748 2804 15804
rect 2804 15748 2808 15804
rect 2744 15744 2808 15748
rect 2824 15804 2888 15808
rect 2824 15748 2828 15804
rect 2828 15748 2884 15804
rect 2884 15748 2888 15804
rect 2824 15744 2888 15748
rect 5847 15804 5911 15808
rect 5847 15748 5851 15804
rect 5851 15748 5907 15804
rect 5907 15748 5911 15804
rect 5847 15744 5911 15748
rect 5927 15804 5991 15808
rect 5927 15748 5931 15804
rect 5931 15748 5987 15804
rect 5987 15748 5991 15804
rect 5927 15744 5991 15748
rect 6007 15804 6071 15808
rect 6007 15748 6011 15804
rect 6011 15748 6067 15804
rect 6067 15748 6071 15804
rect 6007 15744 6071 15748
rect 6087 15804 6151 15808
rect 6087 15748 6091 15804
rect 6091 15748 6147 15804
rect 6147 15748 6151 15804
rect 6087 15744 6151 15748
rect 9111 15804 9175 15808
rect 9111 15748 9115 15804
rect 9115 15748 9171 15804
rect 9171 15748 9175 15804
rect 9111 15744 9175 15748
rect 9191 15804 9255 15808
rect 9191 15748 9195 15804
rect 9195 15748 9251 15804
rect 9251 15748 9255 15804
rect 9191 15744 9255 15748
rect 9271 15804 9335 15808
rect 9271 15748 9275 15804
rect 9275 15748 9331 15804
rect 9331 15748 9335 15804
rect 9271 15744 9335 15748
rect 9351 15804 9415 15808
rect 9351 15748 9355 15804
rect 9355 15748 9411 15804
rect 9411 15748 9415 15804
rect 9351 15744 9415 15748
rect 4215 15260 4279 15264
rect 4215 15204 4219 15260
rect 4219 15204 4275 15260
rect 4275 15204 4279 15260
rect 4215 15200 4279 15204
rect 4295 15260 4359 15264
rect 4295 15204 4299 15260
rect 4299 15204 4355 15260
rect 4355 15204 4359 15260
rect 4295 15200 4359 15204
rect 4375 15260 4439 15264
rect 4375 15204 4379 15260
rect 4379 15204 4435 15260
rect 4435 15204 4439 15260
rect 4375 15200 4439 15204
rect 4455 15260 4519 15264
rect 4455 15204 4459 15260
rect 4459 15204 4515 15260
rect 4515 15204 4519 15260
rect 4455 15200 4519 15204
rect 7479 15260 7543 15264
rect 7479 15204 7483 15260
rect 7483 15204 7539 15260
rect 7539 15204 7543 15260
rect 7479 15200 7543 15204
rect 7559 15260 7623 15264
rect 7559 15204 7563 15260
rect 7563 15204 7619 15260
rect 7619 15204 7623 15260
rect 7559 15200 7623 15204
rect 7639 15260 7703 15264
rect 7639 15204 7643 15260
rect 7643 15204 7699 15260
rect 7699 15204 7703 15260
rect 7639 15200 7703 15204
rect 7719 15260 7783 15264
rect 7719 15204 7723 15260
rect 7723 15204 7779 15260
rect 7779 15204 7783 15260
rect 7719 15200 7783 15204
rect 2584 14716 2648 14720
rect 2584 14660 2588 14716
rect 2588 14660 2644 14716
rect 2644 14660 2648 14716
rect 2584 14656 2648 14660
rect 2664 14716 2728 14720
rect 2664 14660 2668 14716
rect 2668 14660 2724 14716
rect 2724 14660 2728 14716
rect 2664 14656 2728 14660
rect 2744 14716 2808 14720
rect 2744 14660 2748 14716
rect 2748 14660 2804 14716
rect 2804 14660 2808 14716
rect 2744 14656 2808 14660
rect 2824 14716 2888 14720
rect 2824 14660 2828 14716
rect 2828 14660 2884 14716
rect 2884 14660 2888 14716
rect 2824 14656 2888 14660
rect 5847 14716 5911 14720
rect 5847 14660 5851 14716
rect 5851 14660 5907 14716
rect 5907 14660 5911 14716
rect 5847 14656 5911 14660
rect 5927 14716 5991 14720
rect 5927 14660 5931 14716
rect 5931 14660 5987 14716
rect 5987 14660 5991 14716
rect 5927 14656 5991 14660
rect 6007 14716 6071 14720
rect 6007 14660 6011 14716
rect 6011 14660 6067 14716
rect 6067 14660 6071 14716
rect 6007 14656 6071 14660
rect 6087 14716 6151 14720
rect 6087 14660 6091 14716
rect 6091 14660 6147 14716
rect 6147 14660 6151 14716
rect 6087 14656 6151 14660
rect 9111 14716 9175 14720
rect 9111 14660 9115 14716
rect 9115 14660 9171 14716
rect 9171 14660 9175 14716
rect 9111 14656 9175 14660
rect 9191 14716 9255 14720
rect 9191 14660 9195 14716
rect 9195 14660 9251 14716
rect 9251 14660 9255 14716
rect 9191 14656 9255 14660
rect 9271 14716 9335 14720
rect 9271 14660 9275 14716
rect 9275 14660 9331 14716
rect 9331 14660 9335 14716
rect 9271 14656 9335 14660
rect 9351 14716 9415 14720
rect 9351 14660 9355 14716
rect 9355 14660 9411 14716
rect 9411 14660 9415 14716
rect 9351 14656 9415 14660
rect 4215 14172 4279 14176
rect 4215 14116 4219 14172
rect 4219 14116 4275 14172
rect 4275 14116 4279 14172
rect 4215 14112 4279 14116
rect 4295 14172 4359 14176
rect 4295 14116 4299 14172
rect 4299 14116 4355 14172
rect 4355 14116 4359 14172
rect 4295 14112 4359 14116
rect 4375 14172 4439 14176
rect 4375 14116 4379 14172
rect 4379 14116 4435 14172
rect 4435 14116 4439 14172
rect 4375 14112 4439 14116
rect 4455 14172 4519 14176
rect 4455 14116 4459 14172
rect 4459 14116 4515 14172
rect 4515 14116 4519 14172
rect 4455 14112 4519 14116
rect 7479 14172 7543 14176
rect 7479 14116 7483 14172
rect 7483 14116 7539 14172
rect 7539 14116 7543 14172
rect 7479 14112 7543 14116
rect 7559 14172 7623 14176
rect 7559 14116 7563 14172
rect 7563 14116 7619 14172
rect 7619 14116 7623 14172
rect 7559 14112 7623 14116
rect 7639 14172 7703 14176
rect 7639 14116 7643 14172
rect 7643 14116 7699 14172
rect 7699 14116 7703 14172
rect 7639 14112 7703 14116
rect 7719 14172 7783 14176
rect 7719 14116 7723 14172
rect 7723 14116 7779 14172
rect 7779 14116 7783 14172
rect 7719 14112 7783 14116
rect 2584 13628 2648 13632
rect 2584 13572 2588 13628
rect 2588 13572 2644 13628
rect 2644 13572 2648 13628
rect 2584 13568 2648 13572
rect 2664 13628 2728 13632
rect 2664 13572 2668 13628
rect 2668 13572 2724 13628
rect 2724 13572 2728 13628
rect 2664 13568 2728 13572
rect 2744 13628 2808 13632
rect 2744 13572 2748 13628
rect 2748 13572 2804 13628
rect 2804 13572 2808 13628
rect 2744 13568 2808 13572
rect 2824 13628 2888 13632
rect 2824 13572 2828 13628
rect 2828 13572 2884 13628
rect 2884 13572 2888 13628
rect 2824 13568 2888 13572
rect 5847 13628 5911 13632
rect 5847 13572 5851 13628
rect 5851 13572 5907 13628
rect 5907 13572 5911 13628
rect 5847 13568 5911 13572
rect 5927 13628 5991 13632
rect 5927 13572 5931 13628
rect 5931 13572 5987 13628
rect 5987 13572 5991 13628
rect 5927 13568 5991 13572
rect 6007 13628 6071 13632
rect 6007 13572 6011 13628
rect 6011 13572 6067 13628
rect 6067 13572 6071 13628
rect 6007 13568 6071 13572
rect 6087 13628 6151 13632
rect 6087 13572 6091 13628
rect 6091 13572 6147 13628
rect 6147 13572 6151 13628
rect 6087 13568 6151 13572
rect 9111 13628 9175 13632
rect 9111 13572 9115 13628
rect 9115 13572 9171 13628
rect 9171 13572 9175 13628
rect 9111 13568 9175 13572
rect 9191 13628 9255 13632
rect 9191 13572 9195 13628
rect 9195 13572 9251 13628
rect 9251 13572 9255 13628
rect 9191 13568 9255 13572
rect 9271 13628 9335 13632
rect 9271 13572 9275 13628
rect 9275 13572 9331 13628
rect 9331 13572 9335 13628
rect 9271 13568 9335 13572
rect 9351 13628 9415 13632
rect 9351 13572 9355 13628
rect 9355 13572 9411 13628
rect 9411 13572 9415 13628
rect 9351 13568 9415 13572
rect 4215 13084 4279 13088
rect 4215 13028 4219 13084
rect 4219 13028 4275 13084
rect 4275 13028 4279 13084
rect 4215 13024 4279 13028
rect 4295 13084 4359 13088
rect 4295 13028 4299 13084
rect 4299 13028 4355 13084
rect 4355 13028 4359 13084
rect 4295 13024 4359 13028
rect 4375 13084 4439 13088
rect 4375 13028 4379 13084
rect 4379 13028 4435 13084
rect 4435 13028 4439 13084
rect 4375 13024 4439 13028
rect 4455 13084 4519 13088
rect 4455 13028 4459 13084
rect 4459 13028 4515 13084
rect 4515 13028 4519 13084
rect 4455 13024 4519 13028
rect 7479 13084 7543 13088
rect 7479 13028 7483 13084
rect 7483 13028 7539 13084
rect 7539 13028 7543 13084
rect 7479 13024 7543 13028
rect 7559 13084 7623 13088
rect 7559 13028 7563 13084
rect 7563 13028 7619 13084
rect 7619 13028 7623 13084
rect 7559 13024 7623 13028
rect 7639 13084 7703 13088
rect 7639 13028 7643 13084
rect 7643 13028 7699 13084
rect 7699 13028 7703 13084
rect 7639 13024 7703 13028
rect 7719 13084 7783 13088
rect 7719 13028 7723 13084
rect 7723 13028 7779 13084
rect 7779 13028 7783 13084
rect 7719 13024 7783 13028
rect 2584 12540 2648 12544
rect 2584 12484 2588 12540
rect 2588 12484 2644 12540
rect 2644 12484 2648 12540
rect 2584 12480 2648 12484
rect 2664 12540 2728 12544
rect 2664 12484 2668 12540
rect 2668 12484 2724 12540
rect 2724 12484 2728 12540
rect 2664 12480 2728 12484
rect 2744 12540 2808 12544
rect 2744 12484 2748 12540
rect 2748 12484 2804 12540
rect 2804 12484 2808 12540
rect 2744 12480 2808 12484
rect 2824 12540 2888 12544
rect 2824 12484 2828 12540
rect 2828 12484 2884 12540
rect 2884 12484 2888 12540
rect 2824 12480 2888 12484
rect 5847 12540 5911 12544
rect 5847 12484 5851 12540
rect 5851 12484 5907 12540
rect 5907 12484 5911 12540
rect 5847 12480 5911 12484
rect 5927 12540 5991 12544
rect 5927 12484 5931 12540
rect 5931 12484 5987 12540
rect 5987 12484 5991 12540
rect 5927 12480 5991 12484
rect 6007 12540 6071 12544
rect 6007 12484 6011 12540
rect 6011 12484 6067 12540
rect 6067 12484 6071 12540
rect 6007 12480 6071 12484
rect 6087 12540 6151 12544
rect 6087 12484 6091 12540
rect 6091 12484 6147 12540
rect 6147 12484 6151 12540
rect 6087 12480 6151 12484
rect 9111 12540 9175 12544
rect 9111 12484 9115 12540
rect 9115 12484 9171 12540
rect 9171 12484 9175 12540
rect 9111 12480 9175 12484
rect 9191 12540 9255 12544
rect 9191 12484 9195 12540
rect 9195 12484 9251 12540
rect 9251 12484 9255 12540
rect 9191 12480 9255 12484
rect 9271 12540 9335 12544
rect 9271 12484 9275 12540
rect 9275 12484 9331 12540
rect 9331 12484 9335 12540
rect 9271 12480 9335 12484
rect 9351 12540 9415 12544
rect 9351 12484 9355 12540
rect 9355 12484 9411 12540
rect 9411 12484 9415 12540
rect 9351 12480 9415 12484
rect 4215 11996 4279 12000
rect 4215 11940 4219 11996
rect 4219 11940 4275 11996
rect 4275 11940 4279 11996
rect 4215 11936 4279 11940
rect 4295 11996 4359 12000
rect 4295 11940 4299 11996
rect 4299 11940 4355 11996
rect 4355 11940 4359 11996
rect 4295 11936 4359 11940
rect 4375 11996 4439 12000
rect 4375 11940 4379 11996
rect 4379 11940 4435 11996
rect 4435 11940 4439 11996
rect 4375 11936 4439 11940
rect 4455 11996 4519 12000
rect 4455 11940 4459 11996
rect 4459 11940 4515 11996
rect 4515 11940 4519 11996
rect 4455 11936 4519 11940
rect 7479 11996 7543 12000
rect 7479 11940 7483 11996
rect 7483 11940 7539 11996
rect 7539 11940 7543 11996
rect 7479 11936 7543 11940
rect 7559 11996 7623 12000
rect 7559 11940 7563 11996
rect 7563 11940 7619 11996
rect 7619 11940 7623 11996
rect 7559 11936 7623 11940
rect 7639 11996 7703 12000
rect 7639 11940 7643 11996
rect 7643 11940 7699 11996
rect 7699 11940 7703 11996
rect 7639 11936 7703 11940
rect 7719 11996 7783 12000
rect 7719 11940 7723 11996
rect 7723 11940 7779 11996
rect 7779 11940 7783 11996
rect 7719 11936 7783 11940
rect 2584 11452 2648 11456
rect 2584 11396 2588 11452
rect 2588 11396 2644 11452
rect 2644 11396 2648 11452
rect 2584 11392 2648 11396
rect 2664 11452 2728 11456
rect 2664 11396 2668 11452
rect 2668 11396 2724 11452
rect 2724 11396 2728 11452
rect 2664 11392 2728 11396
rect 2744 11452 2808 11456
rect 2744 11396 2748 11452
rect 2748 11396 2804 11452
rect 2804 11396 2808 11452
rect 2744 11392 2808 11396
rect 2824 11452 2888 11456
rect 2824 11396 2828 11452
rect 2828 11396 2884 11452
rect 2884 11396 2888 11452
rect 2824 11392 2888 11396
rect 5847 11452 5911 11456
rect 5847 11396 5851 11452
rect 5851 11396 5907 11452
rect 5907 11396 5911 11452
rect 5847 11392 5911 11396
rect 5927 11452 5991 11456
rect 5927 11396 5931 11452
rect 5931 11396 5987 11452
rect 5987 11396 5991 11452
rect 5927 11392 5991 11396
rect 6007 11452 6071 11456
rect 6007 11396 6011 11452
rect 6011 11396 6067 11452
rect 6067 11396 6071 11452
rect 6007 11392 6071 11396
rect 6087 11452 6151 11456
rect 6087 11396 6091 11452
rect 6091 11396 6147 11452
rect 6147 11396 6151 11452
rect 6087 11392 6151 11396
rect 9111 11452 9175 11456
rect 9111 11396 9115 11452
rect 9115 11396 9171 11452
rect 9171 11396 9175 11452
rect 9111 11392 9175 11396
rect 9191 11452 9255 11456
rect 9191 11396 9195 11452
rect 9195 11396 9251 11452
rect 9251 11396 9255 11452
rect 9191 11392 9255 11396
rect 9271 11452 9335 11456
rect 9271 11396 9275 11452
rect 9275 11396 9331 11452
rect 9331 11396 9335 11452
rect 9271 11392 9335 11396
rect 9351 11452 9415 11456
rect 9351 11396 9355 11452
rect 9355 11396 9411 11452
rect 9411 11396 9415 11452
rect 9351 11392 9415 11396
rect 4215 10908 4279 10912
rect 4215 10852 4219 10908
rect 4219 10852 4275 10908
rect 4275 10852 4279 10908
rect 4215 10848 4279 10852
rect 4295 10908 4359 10912
rect 4295 10852 4299 10908
rect 4299 10852 4355 10908
rect 4355 10852 4359 10908
rect 4295 10848 4359 10852
rect 4375 10908 4439 10912
rect 4375 10852 4379 10908
rect 4379 10852 4435 10908
rect 4435 10852 4439 10908
rect 4375 10848 4439 10852
rect 4455 10908 4519 10912
rect 4455 10852 4459 10908
rect 4459 10852 4515 10908
rect 4515 10852 4519 10908
rect 4455 10848 4519 10852
rect 7479 10908 7543 10912
rect 7479 10852 7483 10908
rect 7483 10852 7539 10908
rect 7539 10852 7543 10908
rect 7479 10848 7543 10852
rect 7559 10908 7623 10912
rect 7559 10852 7563 10908
rect 7563 10852 7619 10908
rect 7619 10852 7623 10908
rect 7559 10848 7623 10852
rect 7639 10908 7703 10912
rect 7639 10852 7643 10908
rect 7643 10852 7699 10908
rect 7699 10852 7703 10908
rect 7639 10848 7703 10852
rect 7719 10908 7783 10912
rect 7719 10852 7723 10908
rect 7723 10852 7779 10908
rect 7779 10852 7783 10908
rect 7719 10848 7783 10852
rect 2584 10364 2648 10368
rect 2584 10308 2588 10364
rect 2588 10308 2644 10364
rect 2644 10308 2648 10364
rect 2584 10304 2648 10308
rect 2664 10364 2728 10368
rect 2664 10308 2668 10364
rect 2668 10308 2724 10364
rect 2724 10308 2728 10364
rect 2664 10304 2728 10308
rect 2744 10364 2808 10368
rect 2744 10308 2748 10364
rect 2748 10308 2804 10364
rect 2804 10308 2808 10364
rect 2744 10304 2808 10308
rect 2824 10364 2888 10368
rect 2824 10308 2828 10364
rect 2828 10308 2884 10364
rect 2884 10308 2888 10364
rect 2824 10304 2888 10308
rect 5847 10364 5911 10368
rect 5847 10308 5851 10364
rect 5851 10308 5907 10364
rect 5907 10308 5911 10364
rect 5847 10304 5911 10308
rect 5927 10364 5991 10368
rect 5927 10308 5931 10364
rect 5931 10308 5987 10364
rect 5987 10308 5991 10364
rect 5927 10304 5991 10308
rect 6007 10364 6071 10368
rect 6007 10308 6011 10364
rect 6011 10308 6067 10364
rect 6067 10308 6071 10364
rect 6007 10304 6071 10308
rect 6087 10364 6151 10368
rect 6087 10308 6091 10364
rect 6091 10308 6147 10364
rect 6147 10308 6151 10364
rect 6087 10304 6151 10308
rect 9111 10364 9175 10368
rect 9111 10308 9115 10364
rect 9115 10308 9171 10364
rect 9171 10308 9175 10364
rect 9111 10304 9175 10308
rect 9191 10364 9255 10368
rect 9191 10308 9195 10364
rect 9195 10308 9251 10364
rect 9251 10308 9255 10364
rect 9191 10304 9255 10308
rect 9271 10364 9335 10368
rect 9271 10308 9275 10364
rect 9275 10308 9331 10364
rect 9331 10308 9335 10364
rect 9271 10304 9335 10308
rect 9351 10364 9415 10368
rect 9351 10308 9355 10364
rect 9355 10308 9411 10364
rect 9411 10308 9415 10364
rect 9351 10304 9415 10308
rect 4215 9820 4279 9824
rect 4215 9764 4219 9820
rect 4219 9764 4275 9820
rect 4275 9764 4279 9820
rect 4215 9760 4279 9764
rect 4295 9820 4359 9824
rect 4295 9764 4299 9820
rect 4299 9764 4355 9820
rect 4355 9764 4359 9820
rect 4295 9760 4359 9764
rect 4375 9820 4439 9824
rect 4375 9764 4379 9820
rect 4379 9764 4435 9820
rect 4435 9764 4439 9820
rect 4375 9760 4439 9764
rect 4455 9820 4519 9824
rect 4455 9764 4459 9820
rect 4459 9764 4515 9820
rect 4515 9764 4519 9820
rect 4455 9760 4519 9764
rect 7479 9820 7543 9824
rect 7479 9764 7483 9820
rect 7483 9764 7539 9820
rect 7539 9764 7543 9820
rect 7479 9760 7543 9764
rect 7559 9820 7623 9824
rect 7559 9764 7563 9820
rect 7563 9764 7619 9820
rect 7619 9764 7623 9820
rect 7559 9760 7623 9764
rect 7639 9820 7703 9824
rect 7639 9764 7643 9820
rect 7643 9764 7699 9820
rect 7699 9764 7703 9820
rect 7639 9760 7703 9764
rect 7719 9820 7783 9824
rect 7719 9764 7723 9820
rect 7723 9764 7779 9820
rect 7779 9764 7783 9820
rect 7719 9760 7783 9764
rect 2584 9276 2648 9280
rect 2584 9220 2588 9276
rect 2588 9220 2644 9276
rect 2644 9220 2648 9276
rect 2584 9216 2648 9220
rect 2664 9276 2728 9280
rect 2664 9220 2668 9276
rect 2668 9220 2724 9276
rect 2724 9220 2728 9276
rect 2664 9216 2728 9220
rect 2744 9276 2808 9280
rect 2744 9220 2748 9276
rect 2748 9220 2804 9276
rect 2804 9220 2808 9276
rect 2744 9216 2808 9220
rect 2824 9276 2888 9280
rect 2824 9220 2828 9276
rect 2828 9220 2884 9276
rect 2884 9220 2888 9276
rect 2824 9216 2888 9220
rect 5847 9276 5911 9280
rect 5847 9220 5851 9276
rect 5851 9220 5907 9276
rect 5907 9220 5911 9276
rect 5847 9216 5911 9220
rect 5927 9276 5991 9280
rect 5927 9220 5931 9276
rect 5931 9220 5987 9276
rect 5987 9220 5991 9276
rect 5927 9216 5991 9220
rect 6007 9276 6071 9280
rect 6007 9220 6011 9276
rect 6011 9220 6067 9276
rect 6067 9220 6071 9276
rect 6007 9216 6071 9220
rect 6087 9276 6151 9280
rect 6087 9220 6091 9276
rect 6091 9220 6147 9276
rect 6147 9220 6151 9276
rect 6087 9216 6151 9220
rect 9111 9276 9175 9280
rect 9111 9220 9115 9276
rect 9115 9220 9171 9276
rect 9171 9220 9175 9276
rect 9111 9216 9175 9220
rect 9191 9276 9255 9280
rect 9191 9220 9195 9276
rect 9195 9220 9251 9276
rect 9251 9220 9255 9276
rect 9191 9216 9255 9220
rect 9271 9276 9335 9280
rect 9271 9220 9275 9276
rect 9275 9220 9331 9276
rect 9331 9220 9335 9276
rect 9271 9216 9335 9220
rect 9351 9276 9415 9280
rect 9351 9220 9355 9276
rect 9355 9220 9411 9276
rect 9411 9220 9415 9276
rect 9351 9216 9415 9220
rect 4215 8732 4279 8736
rect 4215 8676 4219 8732
rect 4219 8676 4275 8732
rect 4275 8676 4279 8732
rect 4215 8672 4279 8676
rect 4295 8732 4359 8736
rect 4295 8676 4299 8732
rect 4299 8676 4355 8732
rect 4355 8676 4359 8732
rect 4295 8672 4359 8676
rect 4375 8732 4439 8736
rect 4375 8676 4379 8732
rect 4379 8676 4435 8732
rect 4435 8676 4439 8732
rect 4375 8672 4439 8676
rect 4455 8732 4519 8736
rect 4455 8676 4459 8732
rect 4459 8676 4515 8732
rect 4515 8676 4519 8732
rect 4455 8672 4519 8676
rect 7479 8732 7543 8736
rect 7479 8676 7483 8732
rect 7483 8676 7539 8732
rect 7539 8676 7543 8732
rect 7479 8672 7543 8676
rect 7559 8732 7623 8736
rect 7559 8676 7563 8732
rect 7563 8676 7619 8732
rect 7619 8676 7623 8732
rect 7559 8672 7623 8676
rect 7639 8732 7703 8736
rect 7639 8676 7643 8732
rect 7643 8676 7699 8732
rect 7699 8676 7703 8732
rect 7639 8672 7703 8676
rect 7719 8732 7783 8736
rect 7719 8676 7723 8732
rect 7723 8676 7779 8732
rect 7779 8676 7783 8732
rect 7719 8672 7783 8676
rect 2584 8188 2648 8192
rect 2584 8132 2588 8188
rect 2588 8132 2644 8188
rect 2644 8132 2648 8188
rect 2584 8128 2648 8132
rect 2664 8188 2728 8192
rect 2664 8132 2668 8188
rect 2668 8132 2724 8188
rect 2724 8132 2728 8188
rect 2664 8128 2728 8132
rect 2744 8188 2808 8192
rect 2744 8132 2748 8188
rect 2748 8132 2804 8188
rect 2804 8132 2808 8188
rect 2744 8128 2808 8132
rect 2824 8188 2888 8192
rect 2824 8132 2828 8188
rect 2828 8132 2884 8188
rect 2884 8132 2888 8188
rect 2824 8128 2888 8132
rect 5847 8188 5911 8192
rect 5847 8132 5851 8188
rect 5851 8132 5907 8188
rect 5907 8132 5911 8188
rect 5847 8128 5911 8132
rect 5927 8188 5991 8192
rect 5927 8132 5931 8188
rect 5931 8132 5987 8188
rect 5987 8132 5991 8188
rect 5927 8128 5991 8132
rect 6007 8188 6071 8192
rect 6007 8132 6011 8188
rect 6011 8132 6067 8188
rect 6067 8132 6071 8188
rect 6007 8128 6071 8132
rect 6087 8188 6151 8192
rect 6087 8132 6091 8188
rect 6091 8132 6147 8188
rect 6147 8132 6151 8188
rect 6087 8128 6151 8132
rect 9111 8188 9175 8192
rect 9111 8132 9115 8188
rect 9115 8132 9171 8188
rect 9171 8132 9175 8188
rect 9111 8128 9175 8132
rect 9191 8188 9255 8192
rect 9191 8132 9195 8188
rect 9195 8132 9251 8188
rect 9251 8132 9255 8188
rect 9191 8128 9255 8132
rect 9271 8188 9335 8192
rect 9271 8132 9275 8188
rect 9275 8132 9331 8188
rect 9331 8132 9335 8188
rect 9271 8128 9335 8132
rect 9351 8188 9415 8192
rect 9351 8132 9355 8188
rect 9355 8132 9411 8188
rect 9411 8132 9415 8188
rect 9351 8128 9415 8132
rect 4215 7644 4279 7648
rect 4215 7588 4219 7644
rect 4219 7588 4275 7644
rect 4275 7588 4279 7644
rect 4215 7584 4279 7588
rect 4295 7644 4359 7648
rect 4295 7588 4299 7644
rect 4299 7588 4355 7644
rect 4355 7588 4359 7644
rect 4295 7584 4359 7588
rect 4375 7644 4439 7648
rect 4375 7588 4379 7644
rect 4379 7588 4435 7644
rect 4435 7588 4439 7644
rect 4375 7584 4439 7588
rect 4455 7644 4519 7648
rect 4455 7588 4459 7644
rect 4459 7588 4515 7644
rect 4515 7588 4519 7644
rect 4455 7584 4519 7588
rect 7479 7644 7543 7648
rect 7479 7588 7483 7644
rect 7483 7588 7539 7644
rect 7539 7588 7543 7644
rect 7479 7584 7543 7588
rect 7559 7644 7623 7648
rect 7559 7588 7563 7644
rect 7563 7588 7619 7644
rect 7619 7588 7623 7644
rect 7559 7584 7623 7588
rect 7639 7644 7703 7648
rect 7639 7588 7643 7644
rect 7643 7588 7699 7644
rect 7699 7588 7703 7644
rect 7639 7584 7703 7588
rect 7719 7644 7783 7648
rect 7719 7588 7723 7644
rect 7723 7588 7779 7644
rect 7779 7588 7783 7644
rect 7719 7584 7783 7588
rect 2584 7100 2648 7104
rect 2584 7044 2588 7100
rect 2588 7044 2644 7100
rect 2644 7044 2648 7100
rect 2584 7040 2648 7044
rect 2664 7100 2728 7104
rect 2664 7044 2668 7100
rect 2668 7044 2724 7100
rect 2724 7044 2728 7100
rect 2664 7040 2728 7044
rect 2744 7100 2808 7104
rect 2744 7044 2748 7100
rect 2748 7044 2804 7100
rect 2804 7044 2808 7100
rect 2744 7040 2808 7044
rect 2824 7100 2888 7104
rect 2824 7044 2828 7100
rect 2828 7044 2884 7100
rect 2884 7044 2888 7100
rect 2824 7040 2888 7044
rect 5847 7100 5911 7104
rect 5847 7044 5851 7100
rect 5851 7044 5907 7100
rect 5907 7044 5911 7100
rect 5847 7040 5911 7044
rect 5927 7100 5991 7104
rect 5927 7044 5931 7100
rect 5931 7044 5987 7100
rect 5987 7044 5991 7100
rect 5927 7040 5991 7044
rect 6007 7100 6071 7104
rect 6007 7044 6011 7100
rect 6011 7044 6067 7100
rect 6067 7044 6071 7100
rect 6007 7040 6071 7044
rect 6087 7100 6151 7104
rect 6087 7044 6091 7100
rect 6091 7044 6147 7100
rect 6147 7044 6151 7100
rect 6087 7040 6151 7044
rect 9111 7100 9175 7104
rect 9111 7044 9115 7100
rect 9115 7044 9171 7100
rect 9171 7044 9175 7100
rect 9111 7040 9175 7044
rect 9191 7100 9255 7104
rect 9191 7044 9195 7100
rect 9195 7044 9251 7100
rect 9251 7044 9255 7100
rect 9191 7040 9255 7044
rect 9271 7100 9335 7104
rect 9271 7044 9275 7100
rect 9275 7044 9331 7100
rect 9331 7044 9335 7100
rect 9271 7040 9335 7044
rect 9351 7100 9415 7104
rect 9351 7044 9355 7100
rect 9355 7044 9411 7100
rect 9411 7044 9415 7100
rect 9351 7040 9415 7044
rect 4215 6556 4279 6560
rect 4215 6500 4219 6556
rect 4219 6500 4275 6556
rect 4275 6500 4279 6556
rect 4215 6496 4279 6500
rect 4295 6556 4359 6560
rect 4295 6500 4299 6556
rect 4299 6500 4355 6556
rect 4355 6500 4359 6556
rect 4295 6496 4359 6500
rect 4375 6556 4439 6560
rect 4375 6500 4379 6556
rect 4379 6500 4435 6556
rect 4435 6500 4439 6556
rect 4375 6496 4439 6500
rect 4455 6556 4519 6560
rect 4455 6500 4459 6556
rect 4459 6500 4515 6556
rect 4515 6500 4519 6556
rect 4455 6496 4519 6500
rect 7479 6556 7543 6560
rect 7479 6500 7483 6556
rect 7483 6500 7539 6556
rect 7539 6500 7543 6556
rect 7479 6496 7543 6500
rect 7559 6556 7623 6560
rect 7559 6500 7563 6556
rect 7563 6500 7619 6556
rect 7619 6500 7623 6556
rect 7559 6496 7623 6500
rect 7639 6556 7703 6560
rect 7639 6500 7643 6556
rect 7643 6500 7699 6556
rect 7699 6500 7703 6556
rect 7639 6496 7703 6500
rect 7719 6556 7783 6560
rect 7719 6500 7723 6556
rect 7723 6500 7779 6556
rect 7779 6500 7783 6556
rect 7719 6496 7783 6500
rect 2584 6012 2648 6016
rect 2584 5956 2588 6012
rect 2588 5956 2644 6012
rect 2644 5956 2648 6012
rect 2584 5952 2648 5956
rect 2664 6012 2728 6016
rect 2664 5956 2668 6012
rect 2668 5956 2724 6012
rect 2724 5956 2728 6012
rect 2664 5952 2728 5956
rect 2744 6012 2808 6016
rect 2744 5956 2748 6012
rect 2748 5956 2804 6012
rect 2804 5956 2808 6012
rect 2744 5952 2808 5956
rect 2824 6012 2888 6016
rect 2824 5956 2828 6012
rect 2828 5956 2884 6012
rect 2884 5956 2888 6012
rect 2824 5952 2888 5956
rect 5847 6012 5911 6016
rect 5847 5956 5851 6012
rect 5851 5956 5907 6012
rect 5907 5956 5911 6012
rect 5847 5952 5911 5956
rect 5927 6012 5991 6016
rect 5927 5956 5931 6012
rect 5931 5956 5987 6012
rect 5987 5956 5991 6012
rect 5927 5952 5991 5956
rect 6007 6012 6071 6016
rect 6007 5956 6011 6012
rect 6011 5956 6067 6012
rect 6067 5956 6071 6012
rect 6007 5952 6071 5956
rect 6087 6012 6151 6016
rect 6087 5956 6091 6012
rect 6091 5956 6147 6012
rect 6147 5956 6151 6012
rect 6087 5952 6151 5956
rect 9111 6012 9175 6016
rect 9111 5956 9115 6012
rect 9115 5956 9171 6012
rect 9171 5956 9175 6012
rect 9111 5952 9175 5956
rect 9191 6012 9255 6016
rect 9191 5956 9195 6012
rect 9195 5956 9251 6012
rect 9251 5956 9255 6012
rect 9191 5952 9255 5956
rect 9271 6012 9335 6016
rect 9271 5956 9275 6012
rect 9275 5956 9331 6012
rect 9331 5956 9335 6012
rect 9271 5952 9335 5956
rect 9351 6012 9415 6016
rect 9351 5956 9355 6012
rect 9355 5956 9411 6012
rect 9411 5956 9415 6012
rect 9351 5952 9415 5956
rect 4215 5468 4279 5472
rect 4215 5412 4219 5468
rect 4219 5412 4275 5468
rect 4275 5412 4279 5468
rect 4215 5408 4279 5412
rect 4295 5468 4359 5472
rect 4295 5412 4299 5468
rect 4299 5412 4355 5468
rect 4355 5412 4359 5468
rect 4295 5408 4359 5412
rect 4375 5468 4439 5472
rect 4375 5412 4379 5468
rect 4379 5412 4435 5468
rect 4435 5412 4439 5468
rect 4375 5408 4439 5412
rect 4455 5468 4519 5472
rect 4455 5412 4459 5468
rect 4459 5412 4515 5468
rect 4515 5412 4519 5468
rect 4455 5408 4519 5412
rect 7479 5468 7543 5472
rect 7479 5412 7483 5468
rect 7483 5412 7539 5468
rect 7539 5412 7543 5468
rect 7479 5408 7543 5412
rect 7559 5468 7623 5472
rect 7559 5412 7563 5468
rect 7563 5412 7619 5468
rect 7619 5412 7623 5468
rect 7559 5408 7623 5412
rect 7639 5468 7703 5472
rect 7639 5412 7643 5468
rect 7643 5412 7699 5468
rect 7699 5412 7703 5468
rect 7639 5408 7703 5412
rect 7719 5468 7783 5472
rect 7719 5412 7723 5468
rect 7723 5412 7779 5468
rect 7779 5412 7783 5468
rect 7719 5408 7783 5412
rect 2584 4924 2648 4928
rect 2584 4868 2588 4924
rect 2588 4868 2644 4924
rect 2644 4868 2648 4924
rect 2584 4864 2648 4868
rect 2664 4924 2728 4928
rect 2664 4868 2668 4924
rect 2668 4868 2724 4924
rect 2724 4868 2728 4924
rect 2664 4864 2728 4868
rect 2744 4924 2808 4928
rect 2744 4868 2748 4924
rect 2748 4868 2804 4924
rect 2804 4868 2808 4924
rect 2744 4864 2808 4868
rect 2824 4924 2888 4928
rect 2824 4868 2828 4924
rect 2828 4868 2884 4924
rect 2884 4868 2888 4924
rect 2824 4864 2888 4868
rect 5847 4924 5911 4928
rect 5847 4868 5851 4924
rect 5851 4868 5907 4924
rect 5907 4868 5911 4924
rect 5847 4864 5911 4868
rect 5927 4924 5991 4928
rect 5927 4868 5931 4924
rect 5931 4868 5987 4924
rect 5987 4868 5991 4924
rect 5927 4864 5991 4868
rect 6007 4924 6071 4928
rect 6007 4868 6011 4924
rect 6011 4868 6067 4924
rect 6067 4868 6071 4924
rect 6007 4864 6071 4868
rect 6087 4924 6151 4928
rect 6087 4868 6091 4924
rect 6091 4868 6147 4924
rect 6147 4868 6151 4924
rect 6087 4864 6151 4868
rect 9111 4924 9175 4928
rect 9111 4868 9115 4924
rect 9115 4868 9171 4924
rect 9171 4868 9175 4924
rect 9111 4864 9175 4868
rect 9191 4924 9255 4928
rect 9191 4868 9195 4924
rect 9195 4868 9251 4924
rect 9251 4868 9255 4924
rect 9191 4864 9255 4868
rect 9271 4924 9335 4928
rect 9271 4868 9275 4924
rect 9275 4868 9331 4924
rect 9331 4868 9335 4924
rect 9271 4864 9335 4868
rect 9351 4924 9415 4928
rect 9351 4868 9355 4924
rect 9355 4868 9411 4924
rect 9411 4868 9415 4924
rect 9351 4864 9415 4868
rect 4215 4380 4279 4384
rect 4215 4324 4219 4380
rect 4219 4324 4275 4380
rect 4275 4324 4279 4380
rect 4215 4320 4279 4324
rect 4295 4380 4359 4384
rect 4295 4324 4299 4380
rect 4299 4324 4355 4380
rect 4355 4324 4359 4380
rect 4295 4320 4359 4324
rect 4375 4380 4439 4384
rect 4375 4324 4379 4380
rect 4379 4324 4435 4380
rect 4435 4324 4439 4380
rect 4375 4320 4439 4324
rect 4455 4380 4519 4384
rect 4455 4324 4459 4380
rect 4459 4324 4515 4380
rect 4515 4324 4519 4380
rect 4455 4320 4519 4324
rect 7479 4380 7543 4384
rect 7479 4324 7483 4380
rect 7483 4324 7539 4380
rect 7539 4324 7543 4380
rect 7479 4320 7543 4324
rect 7559 4380 7623 4384
rect 7559 4324 7563 4380
rect 7563 4324 7619 4380
rect 7619 4324 7623 4380
rect 7559 4320 7623 4324
rect 7639 4380 7703 4384
rect 7639 4324 7643 4380
rect 7643 4324 7699 4380
rect 7699 4324 7703 4380
rect 7639 4320 7703 4324
rect 7719 4380 7783 4384
rect 7719 4324 7723 4380
rect 7723 4324 7779 4380
rect 7779 4324 7783 4380
rect 7719 4320 7783 4324
rect 2584 3836 2648 3840
rect 2584 3780 2588 3836
rect 2588 3780 2644 3836
rect 2644 3780 2648 3836
rect 2584 3776 2648 3780
rect 2664 3836 2728 3840
rect 2664 3780 2668 3836
rect 2668 3780 2724 3836
rect 2724 3780 2728 3836
rect 2664 3776 2728 3780
rect 2744 3836 2808 3840
rect 2744 3780 2748 3836
rect 2748 3780 2804 3836
rect 2804 3780 2808 3836
rect 2744 3776 2808 3780
rect 2824 3836 2888 3840
rect 2824 3780 2828 3836
rect 2828 3780 2884 3836
rect 2884 3780 2888 3836
rect 2824 3776 2888 3780
rect 5847 3836 5911 3840
rect 5847 3780 5851 3836
rect 5851 3780 5907 3836
rect 5907 3780 5911 3836
rect 5847 3776 5911 3780
rect 5927 3836 5991 3840
rect 5927 3780 5931 3836
rect 5931 3780 5987 3836
rect 5987 3780 5991 3836
rect 5927 3776 5991 3780
rect 6007 3836 6071 3840
rect 6007 3780 6011 3836
rect 6011 3780 6067 3836
rect 6067 3780 6071 3836
rect 6007 3776 6071 3780
rect 6087 3836 6151 3840
rect 6087 3780 6091 3836
rect 6091 3780 6147 3836
rect 6147 3780 6151 3836
rect 6087 3776 6151 3780
rect 9111 3836 9175 3840
rect 9111 3780 9115 3836
rect 9115 3780 9171 3836
rect 9171 3780 9175 3836
rect 9111 3776 9175 3780
rect 9191 3836 9255 3840
rect 9191 3780 9195 3836
rect 9195 3780 9251 3836
rect 9251 3780 9255 3836
rect 9191 3776 9255 3780
rect 9271 3836 9335 3840
rect 9271 3780 9275 3836
rect 9275 3780 9331 3836
rect 9331 3780 9335 3836
rect 9271 3776 9335 3780
rect 9351 3836 9415 3840
rect 9351 3780 9355 3836
rect 9355 3780 9411 3836
rect 9411 3780 9415 3836
rect 9351 3776 9415 3780
rect 4215 3292 4279 3296
rect 4215 3236 4219 3292
rect 4219 3236 4275 3292
rect 4275 3236 4279 3292
rect 4215 3232 4279 3236
rect 4295 3292 4359 3296
rect 4295 3236 4299 3292
rect 4299 3236 4355 3292
rect 4355 3236 4359 3292
rect 4295 3232 4359 3236
rect 4375 3292 4439 3296
rect 4375 3236 4379 3292
rect 4379 3236 4435 3292
rect 4435 3236 4439 3292
rect 4375 3232 4439 3236
rect 4455 3292 4519 3296
rect 4455 3236 4459 3292
rect 4459 3236 4515 3292
rect 4515 3236 4519 3292
rect 4455 3232 4519 3236
rect 7479 3292 7543 3296
rect 7479 3236 7483 3292
rect 7483 3236 7539 3292
rect 7539 3236 7543 3292
rect 7479 3232 7543 3236
rect 7559 3292 7623 3296
rect 7559 3236 7563 3292
rect 7563 3236 7619 3292
rect 7619 3236 7623 3292
rect 7559 3232 7623 3236
rect 7639 3292 7703 3296
rect 7639 3236 7643 3292
rect 7643 3236 7699 3292
rect 7699 3236 7703 3292
rect 7639 3232 7703 3236
rect 7719 3292 7783 3296
rect 7719 3236 7723 3292
rect 7723 3236 7779 3292
rect 7779 3236 7783 3292
rect 7719 3232 7783 3236
rect 2584 2748 2648 2752
rect 2584 2692 2588 2748
rect 2588 2692 2644 2748
rect 2644 2692 2648 2748
rect 2584 2688 2648 2692
rect 2664 2748 2728 2752
rect 2664 2692 2668 2748
rect 2668 2692 2724 2748
rect 2724 2692 2728 2748
rect 2664 2688 2728 2692
rect 2744 2748 2808 2752
rect 2744 2692 2748 2748
rect 2748 2692 2804 2748
rect 2804 2692 2808 2748
rect 2744 2688 2808 2692
rect 2824 2748 2888 2752
rect 2824 2692 2828 2748
rect 2828 2692 2884 2748
rect 2884 2692 2888 2748
rect 2824 2688 2888 2692
rect 5847 2748 5911 2752
rect 5847 2692 5851 2748
rect 5851 2692 5907 2748
rect 5907 2692 5911 2748
rect 5847 2688 5911 2692
rect 5927 2748 5991 2752
rect 5927 2692 5931 2748
rect 5931 2692 5987 2748
rect 5987 2692 5991 2748
rect 5927 2688 5991 2692
rect 6007 2748 6071 2752
rect 6007 2692 6011 2748
rect 6011 2692 6067 2748
rect 6067 2692 6071 2748
rect 6007 2688 6071 2692
rect 6087 2748 6151 2752
rect 6087 2692 6091 2748
rect 6091 2692 6147 2748
rect 6147 2692 6151 2748
rect 6087 2688 6151 2692
rect 9111 2748 9175 2752
rect 9111 2692 9115 2748
rect 9115 2692 9171 2748
rect 9171 2692 9175 2748
rect 9111 2688 9175 2692
rect 9191 2748 9255 2752
rect 9191 2692 9195 2748
rect 9195 2692 9251 2748
rect 9251 2692 9255 2748
rect 9191 2688 9255 2692
rect 9271 2748 9335 2752
rect 9271 2692 9275 2748
rect 9275 2692 9331 2748
rect 9331 2692 9335 2748
rect 9271 2688 9335 2692
rect 9351 2748 9415 2752
rect 9351 2692 9355 2748
rect 9355 2692 9411 2748
rect 9411 2692 9415 2748
rect 9351 2688 9415 2692
rect 4215 2204 4279 2208
rect 4215 2148 4219 2204
rect 4219 2148 4275 2204
rect 4275 2148 4279 2204
rect 4215 2144 4279 2148
rect 4295 2204 4359 2208
rect 4295 2148 4299 2204
rect 4299 2148 4355 2204
rect 4355 2148 4359 2204
rect 4295 2144 4359 2148
rect 4375 2204 4439 2208
rect 4375 2148 4379 2204
rect 4379 2148 4435 2204
rect 4435 2148 4439 2204
rect 4375 2144 4439 2148
rect 4455 2204 4519 2208
rect 4455 2148 4459 2204
rect 4459 2148 4515 2204
rect 4515 2148 4519 2204
rect 4455 2144 4519 2148
rect 7479 2204 7543 2208
rect 7479 2148 7483 2204
rect 7483 2148 7539 2204
rect 7539 2148 7543 2204
rect 7479 2144 7543 2148
rect 7559 2204 7623 2208
rect 7559 2148 7563 2204
rect 7563 2148 7619 2204
rect 7619 2148 7623 2204
rect 7559 2144 7623 2148
rect 7639 2204 7703 2208
rect 7639 2148 7643 2204
rect 7643 2148 7699 2204
rect 7699 2148 7703 2204
rect 7639 2144 7703 2148
rect 7719 2204 7783 2208
rect 7719 2148 7723 2204
rect 7723 2148 7779 2204
rect 7779 2148 7783 2204
rect 7719 2144 7783 2148
<< metal4 >>
rect 2575 77824 2896 77840
rect 2575 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2575 76736 2896 77760
rect 2575 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2575 75648 2896 76672
rect 2575 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2575 74560 2896 75584
rect 2575 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2575 73472 2896 74496
rect 2575 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2575 72384 2896 73408
rect 2575 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2575 71296 2896 72320
rect 2575 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2575 70208 2896 71232
rect 2575 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2575 69120 2896 70144
rect 2575 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2575 68032 2896 69056
rect 2575 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2575 66944 2896 67968
rect 2575 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2575 65856 2896 66880
rect 2575 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2575 64768 2896 65792
rect 2575 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2575 63680 2896 64704
rect 2575 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2575 62592 2896 63616
rect 2575 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2575 61504 2896 62528
rect 2575 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2575 60416 2896 61440
rect 2575 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 1715 59396 1781 59397
rect 1715 59332 1716 59396
rect 1780 59332 1781 59396
rect 1715 59331 1781 59332
rect 1718 50965 1778 59331
rect 2575 59328 2896 60352
rect 2575 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2575 58240 2896 59264
rect 2575 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2575 57152 2896 58176
rect 2575 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2575 56064 2896 57088
rect 2575 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2575 54976 2896 56000
rect 2575 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2575 53888 2896 54912
rect 2575 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2575 52800 2896 53824
rect 2575 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2575 51712 2896 52736
rect 2575 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 1715 50964 1781 50965
rect 1715 50900 1716 50964
rect 1780 50900 1781 50964
rect 1715 50899 1781 50900
rect 2575 50624 2896 51648
rect 2575 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2575 49536 2896 50560
rect 2575 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2575 48448 2896 49472
rect 2575 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2575 47360 2896 48384
rect 2575 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2575 46272 2896 47296
rect 4207 77280 4527 77840
rect 4207 77216 4215 77280
rect 4279 77216 4295 77280
rect 4359 77216 4375 77280
rect 4439 77216 4455 77280
rect 4519 77216 4527 77280
rect 4207 76192 4527 77216
rect 4207 76128 4215 76192
rect 4279 76128 4295 76192
rect 4359 76128 4375 76192
rect 4439 76128 4455 76192
rect 4519 76128 4527 76192
rect 4207 75104 4527 76128
rect 4207 75040 4215 75104
rect 4279 75040 4295 75104
rect 4359 75040 4375 75104
rect 4439 75040 4455 75104
rect 4519 75040 4527 75104
rect 4207 74016 4527 75040
rect 4207 73952 4215 74016
rect 4279 73952 4295 74016
rect 4359 73952 4375 74016
rect 4439 73952 4455 74016
rect 4519 73952 4527 74016
rect 4207 72928 4527 73952
rect 4207 72864 4215 72928
rect 4279 72864 4295 72928
rect 4359 72864 4375 72928
rect 4439 72864 4455 72928
rect 4519 72864 4527 72928
rect 4207 71840 4527 72864
rect 4207 71776 4215 71840
rect 4279 71776 4295 71840
rect 4359 71776 4375 71840
rect 4439 71776 4455 71840
rect 4519 71776 4527 71840
rect 4207 70752 4527 71776
rect 4207 70688 4215 70752
rect 4279 70688 4295 70752
rect 4359 70688 4375 70752
rect 4439 70688 4455 70752
rect 4519 70688 4527 70752
rect 4207 69664 4527 70688
rect 4207 69600 4215 69664
rect 4279 69600 4295 69664
rect 4359 69600 4375 69664
rect 4439 69600 4455 69664
rect 4519 69600 4527 69664
rect 4207 68576 4527 69600
rect 4207 68512 4215 68576
rect 4279 68512 4295 68576
rect 4359 68512 4375 68576
rect 4439 68512 4455 68576
rect 4519 68512 4527 68576
rect 4207 67488 4527 68512
rect 4207 67424 4215 67488
rect 4279 67424 4295 67488
rect 4359 67424 4375 67488
rect 4439 67424 4455 67488
rect 4519 67424 4527 67488
rect 4207 66400 4527 67424
rect 4207 66336 4215 66400
rect 4279 66336 4295 66400
rect 4359 66336 4375 66400
rect 4439 66336 4455 66400
rect 4519 66336 4527 66400
rect 4207 65312 4527 66336
rect 4207 65248 4215 65312
rect 4279 65248 4295 65312
rect 4359 65248 4375 65312
rect 4439 65248 4455 65312
rect 4519 65248 4527 65312
rect 4207 64224 4527 65248
rect 4207 64160 4215 64224
rect 4279 64160 4295 64224
rect 4359 64160 4375 64224
rect 4439 64160 4455 64224
rect 4519 64160 4527 64224
rect 4207 63136 4527 64160
rect 4207 63072 4215 63136
rect 4279 63072 4295 63136
rect 4359 63072 4375 63136
rect 4439 63072 4455 63136
rect 4519 63072 4527 63136
rect 4207 62048 4527 63072
rect 4207 61984 4215 62048
rect 4279 61984 4295 62048
rect 4359 61984 4375 62048
rect 4439 61984 4455 62048
rect 4519 61984 4527 62048
rect 4207 60960 4527 61984
rect 4207 60896 4215 60960
rect 4279 60896 4295 60960
rect 4359 60896 4375 60960
rect 4439 60896 4455 60960
rect 4519 60896 4527 60960
rect 4207 59872 4527 60896
rect 4207 59808 4215 59872
rect 4279 59808 4295 59872
rect 4359 59808 4375 59872
rect 4439 59808 4455 59872
rect 4519 59808 4527 59872
rect 4207 58784 4527 59808
rect 4207 58720 4215 58784
rect 4279 58720 4295 58784
rect 4359 58720 4375 58784
rect 4439 58720 4455 58784
rect 4519 58720 4527 58784
rect 4207 57696 4527 58720
rect 4207 57632 4215 57696
rect 4279 57632 4295 57696
rect 4359 57632 4375 57696
rect 4439 57632 4455 57696
rect 4519 57632 4527 57696
rect 4207 56608 4527 57632
rect 4207 56544 4215 56608
rect 4279 56544 4295 56608
rect 4359 56544 4375 56608
rect 4439 56544 4455 56608
rect 4519 56544 4527 56608
rect 4207 55520 4527 56544
rect 4207 55456 4215 55520
rect 4279 55456 4295 55520
rect 4359 55456 4375 55520
rect 4439 55456 4455 55520
rect 4519 55456 4527 55520
rect 4207 54432 4527 55456
rect 4207 54368 4215 54432
rect 4279 54368 4295 54432
rect 4359 54368 4375 54432
rect 4439 54368 4455 54432
rect 4519 54368 4527 54432
rect 4207 53344 4527 54368
rect 4207 53280 4215 53344
rect 4279 53280 4295 53344
rect 4359 53280 4375 53344
rect 4439 53280 4455 53344
rect 4519 53280 4527 53344
rect 4207 52256 4527 53280
rect 4207 52192 4215 52256
rect 4279 52192 4295 52256
rect 4359 52192 4375 52256
rect 4439 52192 4455 52256
rect 4519 52192 4527 52256
rect 4207 51168 4527 52192
rect 4207 51104 4215 51168
rect 4279 51104 4295 51168
rect 4359 51104 4375 51168
rect 4439 51104 4455 51168
rect 4519 51104 4527 51168
rect 4207 50080 4527 51104
rect 4207 50016 4215 50080
rect 4279 50016 4295 50080
rect 4359 50016 4375 50080
rect 4439 50016 4455 50080
rect 4519 50016 4527 50080
rect 4207 48992 4527 50016
rect 4207 48928 4215 48992
rect 4279 48928 4295 48992
rect 4359 48928 4375 48992
rect 4439 48928 4455 48992
rect 4519 48928 4527 48992
rect 4207 47904 4527 48928
rect 4207 47840 4215 47904
rect 4279 47840 4295 47904
rect 4359 47840 4375 47904
rect 4439 47840 4455 47904
rect 4519 47840 4527 47904
rect 3923 47156 3989 47157
rect 3923 47092 3924 47156
rect 3988 47092 3989 47156
rect 3923 47091 3989 47092
rect 2575 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2575 45184 2896 46208
rect 2575 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2575 44096 2896 45120
rect 3926 45117 3986 47091
rect 4207 46816 4527 47840
rect 4207 46752 4215 46816
rect 4279 46752 4295 46816
rect 4359 46752 4375 46816
rect 4439 46752 4455 46816
rect 4519 46752 4527 46816
rect 4207 45728 4527 46752
rect 4207 45664 4215 45728
rect 4279 45664 4295 45728
rect 4359 45664 4375 45728
rect 4439 45664 4455 45728
rect 4519 45664 4527 45728
rect 3923 45116 3989 45117
rect 3923 45052 3924 45116
rect 3988 45052 3989 45116
rect 3923 45051 3989 45052
rect 2575 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2575 43008 2896 44032
rect 2575 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2575 41920 2896 42944
rect 2575 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2575 40832 2896 41856
rect 4207 44640 4527 45664
rect 4207 44576 4215 44640
rect 4279 44576 4295 44640
rect 4359 44576 4375 44640
rect 4439 44576 4455 44640
rect 4519 44576 4527 44640
rect 4207 43552 4527 44576
rect 4207 43488 4215 43552
rect 4279 43488 4295 43552
rect 4359 43488 4375 43552
rect 4439 43488 4455 43552
rect 4519 43488 4527 43552
rect 4207 42464 4527 43488
rect 4207 42400 4215 42464
rect 4279 42400 4295 42464
rect 4359 42400 4375 42464
rect 4439 42400 4455 42464
rect 4519 42400 4527 42464
rect 3003 41852 3069 41853
rect 3003 41788 3004 41852
rect 3068 41788 3069 41852
rect 3003 41787 3069 41788
rect 2575 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2575 39744 2896 40768
rect 3006 40085 3066 41787
rect 4207 41376 4527 42400
rect 5839 77824 6159 77840
rect 5839 77760 5847 77824
rect 5911 77760 5927 77824
rect 5991 77760 6007 77824
rect 6071 77760 6087 77824
rect 6151 77760 6159 77824
rect 5839 76736 6159 77760
rect 5839 76672 5847 76736
rect 5911 76672 5927 76736
rect 5991 76672 6007 76736
rect 6071 76672 6087 76736
rect 6151 76672 6159 76736
rect 5839 75648 6159 76672
rect 5839 75584 5847 75648
rect 5911 75584 5927 75648
rect 5991 75584 6007 75648
rect 6071 75584 6087 75648
rect 6151 75584 6159 75648
rect 5839 74560 6159 75584
rect 5839 74496 5847 74560
rect 5911 74496 5927 74560
rect 5991 74496 6007 74560
rect 6071 74496 6087 74560
rect 6151 74496 6159 74560
rect 5839 73472 6159 74496
rect 5839 73408 5847 73472
rect 5911 73408 5927 73472
rect 5991 73408 6007 73472
rect 6071 73408 6087 73472
rect 6151 73408 6159 73472
rect 5839 72384 6159 73408
rect 5839 72320 5847 72384
rect 5911 72320 5927 72384
rect 5991 72320 6007 72384
rect 6071 72320 6087 72384
rect 6151 72320 6159 72384
rect 5839 71296 6159 72320
rect 5839 71232 5847 71296
rect 5911 71232 5927 71296
rect 5991 71232 6007 71296
rect 6071 71232 6087 71296
rect 6151 71232 6159 71296
rect 5839 70208 6159 71232
rect 5839 70144 5847 70208
rect 5911 70144 5927 70208
rect 5991 70144 6007 70208
rect 6071 70144 6087 70208
rect 6151 70144 6159 70208
rect 5839 69120 6159 70144
rect 5839 69056 5847 69120
rect 5911 69056 5927 69120
rect 5991 69056 6007 69120
rect 6071 69056 6087 69120
rect 6151 69056 6159 69120
rect 5839 68032 6159 69056
rect 5839 67968 5847 68032
rect 5911 67968 5927 68032
rect 5991 67968 6007 68032
rect 6071 67968 6087 68032
rect 6151 67968 6159 68032
rect 5839 66944 6159 67968
rect 5839 66880 5847 66944
rect 5911 66880 5927 66944
rect 5991 66880 6007 66944
rect 6071 66880 6087 66944
rect 6151 66880 6159 66944
rect 5839 65856 6159 66880
rect 5839 65792 5847 65856
rect 5911 65792 5927 65856
rect 5991 65792 6007 65856
rect 6071 65792 6087 65856
rect 6151 65792 6159 65856
rect 5839 64768 6159 65792
rect 5839 64704 5847 64768
rect 5911 64704 5927 64768
rect 5991 64704 6007 64768
rect 6071 64704 6087 64768
rect 6151 64704 6159 64768
rect 5839 63680 6159 64704
rect 5839 63616 5847 63680
rect 5911 63616 5927 63680
rect 5991 63616 6007 63680
rect 6071 63616 6087 63680
rect 6151 63616 6159 63680
rect 5839 62592 6159 63616
rect 5839 62528 5847 62592
rect 5911 62528 5927 62592
rect 5991 62528 6007 62592
rect 6071 62528 6087 62592
rect 6151 62528 6159 62592
rect 5839 61504 6159 62528
rect 5839 61440 5847 61504
rect 5911 61440 5927 61504
rect 5991 61440 6007 61504
rect 6071 61440 6087 61504
rect 6151 61440 6159 61504
rect 5839 60416 6159 61440
rect 5839 60352 5847 60416
rect 5911 60352 5927 60416
rect 5991 60352 6007 60416
rect 6071 60352 6087 60416
rect 6151 60352 6159 60416
rect 5839 59328 6159 60352
rect 5839 59264 5847 59328
rect 5911 59264 5927 59328
rect 5991 59264 6007 59328
rect 6071 59264 6087 59328
rect 6151 59264 6159 59328
rect 5839 58240 6159 59264
rect 5839 58176 5847 58240
rect 5911 58176 5927 58240
rect 5991 58176 6007 58240
rect 6071 58176 6087 58240
rect 6151 58176 6159 58240
rect 5839 57152 6159 58176
rect 5839 57088 5847 57152
rect 5911 57088 5927 57152
rect 5991 57088 6007 57152
rect 6071 57088 6087 57152
rect 6151 57088 6159 57152
rect 5839 56064 6159 57088
rect 5839 56000 5847 56064
rect 5911 56000 5927 56064
rect 5991 56000 6007 56064
rect 6071 56000 6087 56064
rect 6151 56000 6159 56064
rect 5839 54976 6159 56000
rect 5839 54912 5847 54976
rect 5911 54912 5927 54976
rect 5991 54912 6007 54976
rect 6071 54912 6087 54976
rect 6151 54912 6159 54976
rect 5839 53888 6159 54912
rect 5839 53824 5847 53888
rect 5911 53824 5927 53888
rect 5991 53824 6007 53888
rect 6071 53824 6087 53888
rect 6151 53824 6159 53888
rect 5839 52800 6159 53824
rect 5839 52736 5847 52800
rect 5911 52736 5927 52800
rect 5991 52736 6007 52800
rect 6071 52736 6087 52800
rect 6151 52736 6159 52800
rect 5839 51712 6159 52736
rect 5839 51648 5847 51712
rect 5911 51648 5927 51712
rect 5991 51648 6007 51712
rect 6071 51648 6087 51712
rect 6151 51648 6159 51712
rect 5839 50624 6159 51648
rect 5839 50560 5847 50624
rect 5911 50560 5927 50624
rect 5991 50560 6007 50624
rect 6071 50560 6087 50624
rect 6151 50560 6159 50624
rect 5839 49536 6159 50560
rect 5839 49472 5847 49536
rect 5911 49472 5927 49536
rect 5991 49472 6007 49536
rect 6071 49472 6087 49536
rect 6151 49472 6159 49536
rect 5839 48448 6159 49472
rect 5839 48384 5847 48448
rect 5911 48384 5927 48448
rect 5991 48384 6007 48448
rect 6071 48384 6087 48448
rect 6151 48384 6159 48448
rect 5839 47360 6159 48384
rect 5839 47296 5847 47360
rect 5911 47296 5927 47360
rect 5991 47296 6007 47360
rect 6071 47296 6087 47360
rect 6151 47296 6159 47360
rect 5839 46272 6159 47296
rect 5839 46208 5847 46272
rect 5911 46208 5927 46272
rect 5991 46208 6007 46272
rect 6071 46208 6087 46272
rect 6151 46208 6159 46272
rect 5839 45184 6159 46208
rect 5839 45120 5847 45184
rect 5911 45120 5927 45184
rect 5991 45120 6007 45184
rect 6071 45120 6087 45184
rect 6151 45120 6159 45184
rect 5839 44096 6159 45120
rect 5839 44032 5847 44096
rect 5911 44032 5927 44096
rect 5991 44032 6007 44096
rect 6071 44032 6087 44096
rect 6151 44032 6159 44096
rect 5839 43008 6159 44032
rect 5839 42944 5847 43008
rect 5911 42944 5927 43008
rect 5991 42944 6007 43008
rect 6071 42944 6087 43008
rect 6151 42944 6159 43008
rect 5839 41920 6159 42944
rect 5839 41856 5847 41920
rect 5911 41856 5927 41920
rect 5991 41856 6007 41920
rect 6071 41856 6087 41920
rect 6151 41856 6159 41920
rect 4659 41580 4725 41581
rect 4659 41516 4660 41580
rect 4724 41516 4725 41580
rect 4659 41515 4725 41516
rect 4207 41312 4215 41376
rect 4279 41312 4295 41376
rect 4359 41312 4375 41376
rect 4439 41312 4455 41376
rect 4519 41312 4527 41376
rect 4207 40288 4527 41312
rect 4207 40224 4215 40288
rect 4279 40224 4295 40288
rect 4359 40224 4375 40288
rect 4439 40224 4455 40288
rect 4519 40224 4527 40288
rect 3003 40084 3069 40085
rect 3003 40020 3004 40084
rect 3068 40020 3069 40084
rect 3003 40019 3069 40020
rect 2575 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2575 38656 2896 39680
rect 2575 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2575 37568 2896 38592
rect 2575 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2575 36480 2896 37504
rect 2575 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2575 35392 2896 36416
rect 2575 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2575 34304 2896 35328
rect 2575 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2575 33216 2896 34240
rect 2575 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2575 32128 2896 33152
rect 2575 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2575 31040 2896 32064
rect 2575 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2575 29952 2896 30976
rect 2575 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2575 28864 2896 29888
rect 2575 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2575 27776 2896 28800
rect 2575 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2575 26688 2896 27712
rect 2575 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2575 25600 2896 26624
rect 2575 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2575 24512 2896 25536
rect 2575 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2575 23424 2896 24448
rect 2575 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2575 22336 2896 23360
rect 2575 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2575 21248 2896 22272
rect 2575 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2575 20160 2896 21184
rect 2575 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2575 19072 2896 20096
rect 2575 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2575 17984 2896 19008
rect 2575 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2575 16896 2896 17920
rect 2575 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2575 15808 2896 16832
rect 2575 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2575 14720 2896 15744
rect 2575 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2575 13632 2896 14656
rect 2575 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2575 12544 2896 13568
rect 2575 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2575 11456 2896 12480
rect 2575 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2575 10368 2896 11392
rect 2575 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2575 9280 2896 10304
rect 2575 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2575 8192 2896 9216
rect 2575 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2575 7104 2896 8128
rect 2575 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2575 6016 2896 7040
rect 2575 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2575 4928 2896 5952
rect 2575 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2575 3840 2896 4864
rect 2575 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2575 2752 2896 3776
rect 2575 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2575 2128 2896 2688
rect 4207 39200 4527 40224
rect 4207 39136 4215 39200
rect 4279 39136 4295 39200
rect 4359 39136 4375 39200
rect 4439 39136 4455 39200
rect 4519 39136 4527 39200
rect 4207 38112 4527 39136
rect 4207 38048 4215 38112
rect 4279 38048 4295 38112
rect 4359 38048 4375 38112
rect 4439 38048 4455 38112
rect 4519 38048 4527 38112
rect 4207 37024 4527 38048
rect 4207 36960 4215 37024
rect 4279 36960 4295 37024
rect 4359 36960 4375 37024
rect 4439 36960 4455 37024
rect 4519 36960 4527 37024
rect 4207 35936 4527 36960
rect 4207 35872 4215 35936
rect 4279 35872 4295 35936
rect 4359 35872 4375 35936
rect 4439 35872 4455 35936
rect 4519 35872 4527 35936
rect 4207 34848 4527 35872
rect 4207 34784 4215 34848
rect 4279 34784 4295 34848
rect 4359 34784 4375 34848
rect 4439 34784 4455 34848
rect 4519 34784 4527 34848
rect 4207 33760 4527 34784
rect 4662 34373 4722 41515
rect 5839 40832 6159 41856
rect 7471 77280 7791 77840
rect 7471 77216 7479 77280
rect 7543 77216 7559 77280
rect 7623 77216 7639 77280
rect 7703 77216 7719 77280
rect 7783 77216 7791 77280
rect 7471 76192 7791 77216
rect 7471 76128 7479 76192
rect 7543 76128 7559 76192
rect 7623 76128 7639 76192
rect 7703 76128 7719 76192
rect 7783 76128 7791 76192
rect 7471 75104 7791 76128
rect 7471 75040 7479 75104
rect 7543 75040 7559 75104
rect 7623 75040 7639 75104
rect 7703 75040 7719 75104
rect 7783 75040 7791 75104
rect 7471 74016 7791 75040
rect 7471 73952 7479 74016
rect 7543 73952 7559 74016
rect 7623 73952 7639 74016
rect 7703 73952 7719 74016
rect 7783 73952 7791 74016
rect 7471 72928 7791 73952
rect 7471 72864 7479 72928
rect 7543 72864 7559 72928
rect 7623 72864 7639 72928
rect 7703 72864 7719 72928
rect 7783 72864 7791 72928
rect 7471 71840 7791 72864
rect 7471 71776 7479 71840
rect 7543 71776 7559 71840
rect 7623 71776 7639 71840
rect 7703 71776 7719 71840
rect 7783 71776 7791 71840
rect 7471 70752 7791 71776
rect 7471 70688 7479 70752
rect 7543 70688 7559 70752
rect 7623 70688 7639 70752
rect 7703 70688 7719 70752
rect 7783 70688 7791 70752
rect 7471 69664 7791 70688
rect 7471 69600 7479 69664
rect 7543 69600 7559 69664
rect 7623 69600 7639 69664
rect 7703 69600 7719 69664
rect 7783 69600 7791 69664
rect 7471 68576 7791 69600
rect 7471 68512 7479 68576
rect 7543 68512 7559 68576
rect 7623 68512 7639 68576
rect 7703 68512 7719 68576
rect 7783 68512 7791 68576
rect 7471 67488 7791 68512
rect 7471 67424 7479 67488
rect 7543 67424 7559 67488
rect 7623 67424 7639 67488
rect 7703 67424 7719 67488
rect 7783 67424 7791 67488
rect 7471 66400 7791 67424
rect 7471 66336 7479 66400
rect 7543 66336 7559 66400
rect 7623 66336 7639 66400
rect 7703 66336 7719 66400
rect 7783 66336 7791 66400
rect 7471 65312 7791 66336
rect 7471 65248 7479 65312
rect 7543 65248 7559 65312
rect 7623 65248 7639 65312
rect 7703 65248 7719 65312
rect 7783 65248 7791 65312
rect 7471 64224 7791 65248
rect 7471 64160 7479 64224
rect 7543 64160 7559 64224
rect 7623 64160 7639 64224
rect 7703 64160 7719 64224
rect 7783 64160 7791 64224
rect 7471 63136 7791 64160
rect 7471 63072 7479 63136
rect 7543 63072 7559 63136
rect 7623 63072 7639 63136
rect 7703 63072 7719 63136
rect 7783 63072 7791 63136
rect 7471 62048 7791 63072
rect 7471 61984 7479 62048
rect 7543 61984 7559 62048
rect 7623 61984 7639 62048
rect 7703 61984 7719 62048
rect 7783 61984 7791 62048
rect 7471 60960 7791 61984
rect 7471 60896 7479 60960
rect 7543 60896 7559 60960
rect 7623 60896 7639 60960
rect 7703 60896 7719 60960
rect 7783 60896 7791 60960
rect 7471 59872 7791 60896
rect 7471 59808 7479 59872
rect 7543 59808 7559 59872
rect 7623 59808 7639 59872
rect 7703 59808 7719 59872
rect 7783 59808 7791 59872
rect 7471 58784 7791 59808
rect 7471 58720 7479 58784
rect 7543 58720 7559 58784
rect 7623 58720 7639 58784
rect 7703 58720 7719 58784
rect 7783 58720 7791 58784
rect 7471 57696 7791 58720
rect 7471 57632 7479 57696
rect 7543 57632 7559 57696
rect 7623 57632 7639 57696
rect 7703 57632 7719 57696
rect 7783 57632 7791 57696
rect 7471 56608 7791 57632
rect 7471 56544 7479 56608
rect 7543 56544 7559 56608
rect 7623 56544 7639 56608
rect 7703 56544 7719 56608
rect 7783 56544 7791 56608
rect 7471 55520 7791 56544
rect 7471 55456 7479 55520
rect 7543 55456 7559 55520
rect 7623 55456 7639 55520
rect 7703 55456 7719 55520
rect 7783 55456 7791 55520
rect 7471 54432 7791 55456
rect 7471 54368 7479 54432
rect 7543 54368 7559 54432
rect 7623 54368 7639 54432
rect 7703 54368 7719 54432
rect 7783 54368 7791 54432
rect 7471 53344 7791 54368
rect 7471 53280 7479 53344
rect 7543 53280 7559 53344
rect 7623 53280 7639 53344
rect 7703 53280 7719 53344
rect 7783 53280 7791 53344
rect 7471 52256 7791 53280
rect 7471 52192 7479 52256
rect 7543 52192 7559 52256
rect 7623 52192 7639 52256
rect 7703 52192 7719 52256
rect 7783 52192 7791 52256
rect 7471 51168 7791 52192
rect 7471 51104 7479 51168
rect 7543 51104 7559 51168
rect 7623 51104 7639 51168
rect 7703 51104 7719 51168
rect 7783 51104 7791 51168
rect 7471 50080 7791 51104
rect 7471 50016 7479 50080
rect 7543 50016 7559 50080
rect 7623 50016 7639 50080
rect 7703 50016 7719 50080
rect 7783 50016 7791 50080
rect 7471 48992 7791 50016
rect 7471 48928 7479 48992
rect 7543 48928 7559 48992
rect 7623 48928 7639 48992
rect 7703 48928 7719 48992
rect 7783 48928 7791 48992
rect 7471 47904 7791 48928
rect 7471 47840 7479 47904
rect 7543 47840 7559 47904
rect 7623 47840 7639 47904
rect 7703 47840 7719 47904
rect 7783 47840 7791 47904
rect 7471 46816 7791 47840
rect 7471 46752 7479 46816
rect 7543 46752 7559 46816
rect 7623 46752 7639 46816
rect 7703 46752 7719 46816
rect 7783 46752 7791 46816
rect 7471 45728 7791 46752
rect 7471 45664 7479 45728
rect 7543 45664 7559 45728
rect 7623 45664 7639 45728
rect 7703 45664 7719 45728
rect 7783 45664 7791 45728
rect 7471 44640 7791 45664
rect 7471 44576 7479 44640
rect 7543 44576 7559 44640
rect 7623 44576 7639 44640
rect 7703 44576 7719 44640
rect 7783 44576 7791 44640
rect 7471 43552 7791 44576
rect 7471 43488 7479 43552
rect 7543 43488 7559 43552
rect 7623 43488 7639 43552
rect 7703 43488 7719 43552
rect 7783 43488 7791 43552
rect 7471 42464 7791 43488
rect 7471 42400 7479 42464
rect 7543 42400 7559 42464
rect 7623 42400 7639 42464
rect 7703 42400 7719 42464
rect 7783 42400 7791 42464
rect 7471 41376 7791 42400
rect 7471 41312 7479 41376
rect 7543 41312 7559 41376
rect 7623 41312 7639 41376
rect 7703 41312 7719 41376
rect 7783 41312 7791 41376
rect 6499 41308 6565 41309
rect 6499 41244 6500 41308
rect 6564 41244 6565 41308
rect 6499 41243 6565 41244
rect 5839 40768 5847 40832
rect 5911 40768 5927 40832
rect 5991 40768 6007 40832
rect 6071 40768 6087 40832
rect 6151 40768 6159 40832
rect 5839 39744 6159 40768
rect 5839 39680 5847 39744
rect 5911 39680 5927 39744
rect 5991 39680 6007 39744
rect 6071 39680 6087 39744
rect 6151 39680 6159 39744
rect 5839 38656 6159 39680
rect 5839 38592 5847 38656
rect 5911 38592 5927 38656
rect 5991 38592 6007 38656
rect 6071 38592 6087 38656
rect 6151 38592 6159 38656
rect 5839 37568 6159 38592
rect 5839 37504 5847 37568
rect 5911 37504 5927 37568
rect 5991 37504 6007 37568
rect 6071 37504 6087 37568
rect 6151 37504 6159 37568
rect 5839 36480 6159 37504
rect 6502 36957 6562 41243
rect 7471 40288 7791 41312
rect 7471 40224 7479 40288
rect 7543 40224 7559 40288
rect 7623 40224 7639 40288
rect 7703 40224 7719 40288
rect 7783 40224 7791 40288
rect 7471 39200 7791 40224
rect 7471 39136 7479 39200
rect 7543 39136 7559 39200
rect 7623 39136 7639 39200
rect 7703 39136 7719 39200
rect 7783 39136 7791 39200
rect 7471 38112 7791 39136
rect 7471 38048 7479 38112
rect 7543 38048 7559 38112
rect 7623 38048 7639 38112
rect 7703 38048 7719 38112
rect 7783 38048 7791 38112
rect 7471 37024 7791 38048
rect 7471 36960 7479 37024
rect 7543 36960 7559 37024
rect 7623 36960 7639 37024
rect 7703 36960 7719 37024
rect 7783 36960 7791 37024
rect 6499 36956 6565 36957
rect 6499 36892 6500 36956
rect 6564 36892 6565 36956
rect 6499 36891 6565 36892
rect 5839 36416 5847 36480
rect 5911 36416 5927 36480
rect 5991 36416 6007 36480
rect 6071 36416 6087 36480
rect 6151 36416 6159 36480
rect 5839 35392 6159 36416
rect 5839 35328 5847 35392
rect 5911 35328 5927 35392
rect 5991 35328 6007 35392
rect 6071 35328 6087 35392
rect 6151 35328 6159 35392
rect 4659 34372 4725 34373
rect 4659 34308 4660 34372
rect 4724 34308 4725 34372
rect 4659 34307 4725 34308
rect 4207 33696 4215 33760
rect 4279 33696 4295 33760
rect 4359 33696 4375 33760
rect 4439 33696 4455 33760
rect 4519 33696 4527 33760
rect 4207 32672 4527 33696
rect 4207 32608 4215 32672
rect 4279 32608 4295 32672
rect 4359 32608 4375 32672
rect 4439 32608 4455 32672
rect 4519 32608 4527 32672
rect 4207 31584 4527 32608
rect 4207 31520 4215 31584
rect 4279 31520 4295 31584
rect 4359 31520 4375 31584
rect 4439 31520 4455 31584
rect 4519 31520 4527 31584
rect 4207 30496 4527 31520
rect 4207 30432 4215 30496
rect 4279 30432 4295 30496
rect 4359 30432 4375 30496
rect 4439 30432 4455 30496
rect 4519 30432 4527 30496
rect 4207 29408 4527 30432
rect 4207 29344 4215 29408
rect 4279 29344 4295 29408
rect 4359 29344 4375 29408
rect 4439 29344 4455 29408
rect 4519 29344 4527 29408
rect 4207 28320 4527 29344
rect 4207 28256 4215 28320
rect 4279 28256 4295 28320
rect 4359 28256 4375 28320
rect 4439 28256 4455 28320
rect 4519 28256 4527 28320
rect 4207 27232 4527 28256
rect 4207 27168 4215 27232
rect 4279 27168 4295 27232
rect 4359 27168 4375 27232
rect 4439 27168 4455 27232
rect 4519 27168 4527 27232
rect 4207 26144 4527 27168
rect 4207 26080 4215 26144
rect 4279 26080 4295 26144
rect 4359 26080 4375 26144
rect 4439 26080 4455 26144
rect 4519 26080 4527 26144
rect 4207 25056 4527 26080
rect 4207 24992 4215 25056
rect 4279 24992 4295 25056
rect 4359 24992 4375 25056
rect 4439 24992 4455 25056
rect 4519 24992 4527 25056
rect 4207 23968 4527 24992
rect 4207 23904 4215 23968
rect 4279 23904 4295 23968
rect 4359 23904 4375 23968
rect 4439 23904 4455 23968
rect 4519 23904 4527 23968
rect 4207 22880 4527 23904
rect 4207 22816 4215 22880
rect 4279 22816 4295 22880
rect 4359 22816 4375 22880
rect 4439 22816 4455 22880
rect 4519 22816 4527 22880
rect 4207 21792 4527 22816
rect 4207 21728 4215 21792
rect 4279 21728 4295 21792
rect 4359 21728 4375 21792
rect 4439 21728 4455 21792
rect 4519 21728 4527 21792
rect 4207 20704 4527 21728
rect 4207 20640 4215 20704
rect 4279 20640 4295 20704
rect 4359 20640 4375 20704
rect 4439 20640 4455 20704
rect 4519 20640 4527 20704
rect 4207 19616 4527 20640
rect 4207 19552 4215 19616
rect 4279 19552 4295 19616
rect 4359 19552 4375 19616
rect 4439 19552 4455 19616
rect 4519 19552 4527 19616
rect 4207 18528 4527 19552
rect 4207 18464 4215 18528
rect 4279 18464 4295 18528
rect 4359 18464 4375 18528
rect 4439 18464 4455 18528
rect 4519 18464 4527 18528
rect 4207 17440 4527 18464
rect 4207 17376 4215 17440
rect 4279 17376 4295 17440
rect 4359 17376 4375 17440
rect 4439 17376 4455 17440
rect 4519 17376 4527 17440
rect 4207 16352 4527 17376
rect 4207 16288 4215 16352
rect 4279 16288 4295 16352
rect 4359 16288 4375 16352
rect 4439 16288 4455 16352
rect 4519 16288 4527 16352
rect 4207 15264 4527 16288
rect 4207 15200 4215 15264
rect 4279 15200 4295 15264
rect 4359 15200 4375 15264
rect 4439 15200 4455 15264
rect 4519 15200 4527 15264
rect 4207 14176 4527 15200
rect 4207 14112 4215 14176
rect 4279 14112 4295 14176
rect 4359 14112 4375 14176
rect 4439 14112 4455 14176
rect 4519 14112 4527 14176
rect 4207 13088 4527 14112
rect 4207 13024 4215 13088
rect 4279 13024 4295 13088
rect 4359 13024 4375 13088
rect 4439 13024 4455 13088
rect 4519 13024 4527 13088
rect 4207 12000 4527 13024
rect 4207 11936 4215 12000
rect 4279 11936 4295 12000
rect 4359 11936 4375 12000
rect 4439 11936 4455 12000
rect 4519 11936 4527 12000
rect 4207 10912 4527 11936
rect 4207 10848 4215 10912
rect 4279 10848 4295 10912
rect 4359 10848 4375 10912
rect 4439 10848 4455 10912
rect 4519 10848 4527 10912
rect 4207 9824 4527 10848
rect 4207 9760 4215 9824
rect 4279 9760 4295 9824
rect 4359 9760 4375 9824
rect 4439 9760 4455 9824
rect 4519 9760 4527 9824
rect 4207 8736 4527 9760
rect 4207 8672 4215 8736
rect 4279 8672 4295 8736
rect 4359 8672 4375 8736
rect 4439 8672 4455 8736
rect 4519 8672 4527 8736
rect 4207 7648 4527 8672
rect 4207 7584 4215 7648
rect 4279 7584 4295 7648
rect 4359 7584 4375 7648
rect 4439 7584 4455 7648
rect 4519 7584 4527 7648
rect 4207 6560 4527 7584
rect 4207 6496 4215 6560
rect 4279 6496 4295 6560
rect 4359 6496 4375 6560
rect 4439 6496 4455 6560
rect 4519 6496 4527 6560
rect 4207 5472 4527 6496
rect 4207 5408 4215 5472
rect 4279 5408 4295 5472
rect 4359 5408 4375 5472
rect 4439 5408 4455 5472
rect 4519 5408 4527 5472
rect 4207 4384 4527 5408
rect 4207 4320 4215 4384
rect 4279 4320 4295 4384
rect 4359 4320 4375 4384
rect 4439 4320 4455 4384
rect 4519 4320 4527 4384
rect 4207 3296 4527 4320
rect 4207 3232 4215 3296
rect 4279 3232 4295 3296
rect 4359 3232 4375 3296
rect 4439 3232 4455 3296
rect 4519 3232 4527 3296
rect 4207 2208 4527 3232
rect 4207 2144 4215 2208
rect 4279 2144 4295 2208
rect 4359 2144 4375 2208
rect 4439 2144 4455 2208
rect 4519 2144 4527 2208
rect 4207 2128 4527 2144
rect 5839 34304 6159 35328
rect 5839 34240 5847 34304
rect 5911 34240 5927 34304
rect 5991 34240 6007 34304
rect 6071 34240 6087 34304
rect 6151 34240 6159 34304
rect 5839 33216 6159 34240
rect 5839 33152 5847 33216
rect 5911 33152 5927 33216
rect 5991 33152 6007 33216
rect 6071 33152 6087 33216
rect 6151 33152 6159 33216
rect 5839 32128 6159 33152
rect 5839 32064 5847 32128
rect 5911 32064 5927 32128
rect 5991 32064 6007 32128
rect 6071 32064 6087 32128
rect 6151 32064 6159 32128
rect 5839 31040 6159 32064
rect 5839 30976 5847 31040
rect 5911 30976 5927 31040
rect 5991 30976 6007 31040
rect 6071 30976 6087 31040
rect 6151 30976 6159 31040
rect 5839 29952 6159 30976
rect 5839 29888 5847 29952
rect 5911 29888 5927 29952
rect 5991 29888 6007 29952
rect 6071 29888 6087 29952
rect 6151 29888 6159 29952
rect 5839 28864 6159 29888
rect 5839 28800 5847 28864
rect 5911 28800 5927 28864
rect 5991 28800 6007 28864
rect 6071 28800 6087 28864
rect 6151 28800 6159 28864
rect 5839 27776 6159 28800
rect 5839 27712 5847 27776
rect 5911 27712 5927 27776
rect 5991 27712 6007 27776
rect 6071 27712 6087 27776
rect 6151 27712 6159 27776
rect 5839 26688 6159 27712
rect 5839 26624 5847 26688
rect 5911 26624 5927 26688
rect 5991 26624 6007 26688
rect 6071 26624 6087 26688
rect 6151 26624 6159 26688
rect 5839 25600 6159 26624
rect 5839 25536 5847 25600
rect 5911 25536 5927 25600
rect 5991 25536 6007 25600
rect 6071 25536 6087 25600
rect 6151 25536 6159 25600
rect 5839 24512 6159 25536
rect 5839 24448 5847 24512
rect 5911 24448 5927 24512
rect 5991 24448 6007 24512
rect 6071 24448 6087 24512
rect 6151 24448 6159 24512
rect 5839 23424 6159 24448
rect 5839 23360 5847 23424
rect 5911 23360 5927 23424
rect 5991 23360 6007 23424
rect 6071 23360 6087 23424
rect 6151 23360 6159 23424
rect 5839 22336 6159 23360
rect 5839 22272 5847 22336
rect 5911 22272 5927 22336
rect 5991 22272 6007 22336
rect 6071 22272 6087 22336
rect 6151 22272 6159 22336
rect 5839 21248 6159 22272
rect 5839 21184 5847 21248
rect 5911 21184 5927 21248
rect 5991 21184 6007 21248
rect 6071 21184 6087 21248
rect 6151 21184 6159 21248
rect 5839 20160 6159 21184
rect 5839 20096 5847 20160
rect 5911 20096 5927 20160
rect 5991 20096 6007 20160
rect 6071 20096 6087 20160
rect 6151 20096 6159 20160
rect 5839 19072 6159 20096
rect 5839 19008 5847 19072
rect 5911 19008 5927 19072
rect 5991 19008 6007 19072
rect 6071 19008 6087 19072
rect 6151 19008 6159 19072
rect 5839 17984 6159 19008
rect 5839 17920 5847 17984
rect 5911 17920 5927 17984
rect 5991 17920 6007 17984
rect 6071 17920 6087 17984
rect 6151 17920 6159 17984
rect 5839 16896 6159 17920
rect 5839 16832 5847 16896
rect 5911 16832 5927 16896
rect 5991 16832 6007 16896
rect 6071 16832 6087 16896
rect 6151 16832 6159 16896
rect 5839 15808 6159 16832
rect 5839 15744 5847 15808
rect 5911 15744 5927 15808
rect 5991 15744 6007 15808
rect 6071 15744 6087 15808
rect 6151 15744 6159 15808
rect 5839 14720 6159 15744
rect 5839 14656 5847 14720
rect 5911 14656 5927 14720
rect 5991 14656 6007 14720
rect 6071 14656 6087 14720
rect 6151 14656 6159 14720
rect 5839 13632 6159 14656
rect 5839 13568 5847 13632
rect 5911 13568 5927 13632
rect 5991 13568 6007 13632
rect 6071 13568 6087 13632
rect 6151 13568 6159 13632
rect 5839 12544 6159 13568
rect 5839 12480 5847 12544
rect 5911 12480 5927 12544
rect 5991 12480 6007 12544
rect 6071 12480 6087 12544
rect 6151 12480 6159 12544
rect 5839 11456 6159 12480
rect 5839 11392 5847 11456
rect 5911 11392 5927 11456
rect 5991 11392 6007 11456
rect 6071 11392 6087 11456
rect 6151 11392 6159 11456
rect 5839 10368 6159 11392
rect 5839 10304 5847 10368
rect 5911 10304 5927 10368
rect 5991 10304 6007 10368
rect 6071 10304 6087 10368
rect 6151 10304 6159 10368
rect 5839 9280 6159 10304
rect 5839 9216 5847 9280
rect 5911 9216 5927 9280
rect 5991 9216 6007 9280
rect 6071 9216 6087 9280
rect 6151 9216 6159 9280
rect 5839 8192 6159 9216
rect 5839 8128 5847 8192
rect 5911 8128 5927 8192
rect 5991 8128 6007 8192
rect 6071 8128 6087 8192
rect 6151 8128 6159 8192
rect 5839 7104 6159 8128
rect 5839 7040 5847 7104
rect 5911 7040 5927 7104
rect 5991 7040 6007 7104
rect 6071 7040 6087 7104
rect 6151 7040 6159 7104
rect 5839 6016 6159 7040
rect 5839 5952 5847 6016
rect 5911 5952 5927 6016
rect 5991 5952 6007 6016
rect 6071 5952 6087 6016
rect 6151 5952 6159 6016
rect 5839 4928 6159 5952
rect 5839 4864 5847 4928
rect 5911 4864 5927 4928
rect 5991 4864 6007 4928
rect 6071 4864 6087 4928
rect 6151 4864 6159 4928
rect 5839 3840 6159 4864
rect 5839 3776 5847 3840
rect 5911 3776 5927 3840
rect 5991 3776 6007 3840
rect 6071 3776 6087 3840
rect 6151 3776 6159 3840
rect 5839 2752 6159 3776
rect 5839 2688 5847 2752
rect 5911 2688 5927 2752
rect 5991 2688 6007 2752
rect 6071 2688 6087 2752
rect 6151 2688 6159 2752
rect 5839 2128 6159 2688
rect 7471 35936 7791 36960
rect 7471 35872 7479 35936
rect 7543 35872 7559 35936
rect 7623 35872 7639 35936
rect 7703 35872 7719 35936
rect 7783 35872 7791 35936
rect 7471 34848 7791 35872
rect 7471 34784 7479 34848
rect 7543 34784 7559 34848
rect 7623 34784 7639 34848
rect 7703 34784 7719 34848
rect 7783 34784 7791 34848
rect 7471 33760 7791 34784
rect 7471 33696 7479 33760
rect 7543 33696 7559 33760
rect 7623 33696 7639 33760
rect 7703 33696 7719 33760
rect 7783 33696 7791 33760
rect 7471 32672 7791 33696
rect 7471 32608 7479 32672
rect 7543 32608 7559 32672
rect 7623 32608 7639 32672
rect 7703 32608 7719 32672
rect 7783 32608 7791 32672
rect 7471 31584 7791 32608
rect 7471 31520 7479 31584
rect 7543 31520 7559 31584
rect 7623 31520 7639 31584
rect 7703 31520 7719 31584
rect 7783 31520 7791 31584
rect 7471 30496 7791 31520
rect 7471 30432 7479 30496
rect 7543 30432 7559 30496
rect 7623 30432 7639 30496
rect 7703 30432 7719 30496
rect 7783 30432 7791 30496
rect 7471 29408 7791 30432
rect 7471 29344 7479 29408
rect 7543 29344 7559 29408
rect 7623 29344 7639 29408
rect 7703 29344 7719 29408
rect 7783 29344 7791 29408
rect 7471 28320 7791 29344
rect 7471 28256 7479 28320
rect 7543 28256 7559 28320
rect 7623 28256 7639 28320
rect 7703 28256 7719 28320
rect 7783 28256 7791 28320
rect 7471 27232 7791 28256
rect 7471 27168 7479 27232
rect 7543 27168 7559 27232
rect 7623 27168 7639 27232
rect 7703 27168 7719 27232
rect 7783 27168 7791 27232
rect 7471 26144 7791 27168
rect 7471 26080 7479 26144
rect 7543 26080 7559 26144
rect 7623 26080 7639 26144
rect 7703 26080 7719 26144
rect 7783 26080 7791 26144
rect 7471 25056 7791 26080
rect 7471 24992 7479 25056
rect 7543 24992 7559 25056
rect 7623 24992 7639 25056
rect 7703 24992 7719 25056
rect 7783 24992 7791 25056
rect 7471 23968 7791 24992
rect 7471 23904 7479 23968
rect 7543 23904 7559 23968
rect 7623 23904 7639 23968
rect 7703 23904 7719 23968
rect 7783 23904 7791 23968
rect 7471 22880 7791 23904
rect 7471 22816 7479 22880
rect 7543 22816 7559 22880
rect 7623 22816 7639 22880
rect 7703 22816 7719 22880
rect 7783 22816 7791 22880
rect 7471 21792 7791 22816
rect 7471 21728 7479 21792
rect 7543 21728 7559 21792
rect 7623 21728 7639 21792
rect 7703 21728 7719 21792
rect 7783 21728 7791 21792
rect 7471 20704 7791 21728
rect 7471 20640 7479 20704
rect 7543 20640 7559 20704
rect 7623 20640 7639 20704
rect 7703 20640 7719 20704
rect 7783 20640 7791 20704
rect 7471 19616 7791 20640
rect 7471 19552 7479 19616
rect 7543 19552 7559 19616
rect 7623 19552 7639 19616
rect 7703 19552 7719 19616
rect 7783 19552 7791 19616
rect 7471 18528 7791 19552
rect 7471 18464 7479 18528
rect 7543 18464 7559 18528
rect 7623 18464 7639 18528
rect 7703 18464 7719 18528
rect 7783 18464 7791 18528
rect 7471 17440 7791 18464
rect 7471 17376 7479 17440
rect 7543 17376 7559 17440
rect 7623 17376 7639 17440
rect 7703 17376 7719 17440
rect 7783 17376 7791 17440
rect 7471 16352 7791 17376
rect 7471 16288 7479 16352
rect 7543 16288 7559 16352
rect 7623 16288 7639 16352
rect 7703 16288 7719 16352
rect 7783 16288 7791 16352
rect 7471 15264 7791 16288
rect 7471 15200 7479 15264
rect 7543 15200 7559 15264
rect 7623 15200 7639 15264
rect 7703 15200 7719 15264
rect 7783 15200 7791 15264
rect 7471 14176 7791 15200
rect 7471 14112 7479 14176
rect 7543 14112 7559 14176
rect 7623 14112 7639 14176
rect 7703 14112 7719 14176
rect 7783 14112 7791 14176
rect 7471 13088 7791 14112
rect 7471 13024 7479 13088
rect 7543 13024 7559 13088
rect 7623 13024 7639 13088
rect 7703 13024 7719 13088
rect 7783 13024 7791 13088
rect 7471 12000 7791 13024
rect 7471 11936 7479 12000
rect 7543 11936 7559 12000
rect 7623 11936 7639 12000
rect 7703 11936 7719 12000
rect 7783 11936 7791 12000
rect 7471 10912 7791 11936
rect 7471 10848 7479 10912
rect 7543 10848 7559 10912
rect 7623 10848 7639 10912
rect 7703 10848 7719 10912
rect 7783 10848 7791 10912
rect 7471 9824 7791 10848
rect 7471 9760 7479 9824
rect 7543 9760 7559 9824
rect 7623 9760 7639 9824
rect 7703 9760 7719 9824
rect 7783 9760 7791 9824
rect 7471 8736 7791 9760
rect 7471 8672 7479 8736
rect 7543 8672 7559 8736
rect 7623 8672 7639 8736
rect 7703 8672 7719 8736
rect 7783 8672 7791 8736
rect 7471 7648 7791 8672
rect 7471 7584 7479 7648
rect 7543 7584 7559 7648
rect 7623 7584 7639 7648
rect 7703 7584 7719 7648
rect 7783 7584 7791 7648
rect 7471 6560 7791 7584
rect 7471 6496 7479 6560
rect 7543 6496 7559 6560
rect 7623 6496 7639 6560
rect 7703 6496 7719 6560
rect 7783 6496 7791 6560
rect 7471 5472 7791 6496
rect 7471 5408 7479 5472
rect 7543 5408 7559 5472
rect 7623 5408 7639 5472
rect 7703 5408 7719 5472
rect 7783 5408 7791 5472
rect 7471 4384 7791 5408
rect 7471 4320 7479 4384
rect 7543 4320 7559 4384
rect 7623 4320 7639 4384
rect 7703 4320 7719 4384
rect 7783 4320 7791 4384
rect 7471 3296 7791 4320
rect 7471 3232 7479 3296
rect 7543 3232 7559 3296
rect 7623 3232 7639 3296
rect 7703 3232 7719 3296
rect 7783 3232 7791 3296
rect 7471 2208 7791 3232
rect 7471 2144 7479 2208
rect 7543 2144 7559 2208
rect 7623 2144 7639 2208
rect 7703 2144 7719 2208
rect 7783 2144 7791 2208
rect 7471 2128 7791 2144
rect 9103 77824 9423 77840
rect 9103 77760 9111 77824
rect 9175 77760 9191 77824
rect 9255 77760 9271 77824
rect 9335 77760 9351 77824
rect 9415 77760 9423 77824
rect 9103 76736 9423 77760
rect 9103 76672 9111 76736
rect 9175 76672 9191 76736
rect 9255 76672 9271 76736
rect 9335 76672 9351 76736
rect 9415 76672 9423 76736
rect 9103 75648 9423 76672
rect 9103 75584 9111 75648
rect 9175 75584 9191 75648
rect 9255 75584 9271 75648
rect 9335 75584 9351 75648
rect 9415 75584 9423 75648
rect 9103 74560 9423 75584
rect 9103 74496 9111 74560
rect 9175 74496 9191 74560
rect 9255 74496 9271 74560
rect 9335 74496 9351 74560
rect 9415 74496 9423 74560
rect 9103 73472 9423 74496
rect 9103 73408 9111 73472
rect 9175 73408 9191 73472
rect 9255 73408 9271 73472
rect 9335 73408 9351 73472
rect 9415 73408 9423 73472
rect 9103 72384 9423 73408
rect 9103 72320 9111 72384
rect 9175 72320 9191 72384
rect 9255 72320 9271 72384
rect 9335 72320 9351 72384
rect 9415 72320 9423 72384
rect 9103 71296 9423 72320
rect 9103 71232 9111 71296
rect 9175 71232 9191 71296
rect 9255 71232 9271 71296
rect 9335 71232 9351 71296
rect 9415 71232 9423 71296
rect 9103 70208 9423 71232
rect 9103 70144 9111 70208
rect 9175 70144 9191 70208
rect 9255 70144 9271 70208
rect 9335 70144 9351 70208
rect 9415 70144 9423 70208
rect 9103 69120 9423 70144
rect 9103 69056 9111 69120
rect 9175 69056 9191 69120
rect 9255 69056 9271 69120
rect 9335 69056 9351 69120
rect 9415 69056 9423 69120
rect 9103 68032 9423 69056
rect 9103 67968 9111 68032
rect 9175 67968 9191 68032
rect 9255 67968 9271 68032
rect 9335 67968 9351 68032
rect 9415 67968 9423 68032
rect 9103 66944 9423 67968
rect 9103 66880 9111 66944
rect 9175 66880 9191 66944
rect 9255 66880 9271 66944
rect 9335 66880 9351 66944
rect 9415 66880 9423 66944
rect 9103 65856 9423 66880
rect 9103 65792 9111 65856
rect 9175 65792 9191 65856
rect 9255 65792 9271 65856
rect 9335 65792 9351 65856
rect 9415 65792 9423 65856
rect 9103 64768 9423 65792
rect 9103 64704 9111 64768
rect 9175 64704 9191 64768
rect 9255 64704 9271 64768
rect 9335 64704 9351 64768
rect 9415 64704 9423 64768
rect 9103 63680 9423 64704
rect 9103 63616 9111 63680
rect 9175 63616 9191 63680
rect 9255 63616 9271 63680
rect 9335 63616 9351 63680
rect 9415 63616 9423 63680
rect 9103 62592 9423 63616
rect 9103 62528 9111 62592
rect 9175 62528 9191 62592
rect 9255 62528 9271 62592
rect 9335 62528 9351 62592
rect 9415 62528 9423 62592
rect 9103 61504 9423 62528
rect 9103 61440 9111 61504
rect 9175 61440 9191 61504
rect 9255 61440 9271 61504
rect 9335 61440 9351 61504
rect 9415 61440 9423 61504
rect 9103 60416 9423 61440
rect 9103 60352 9111 60416
rect 9175 60352 9191 60416
rect 9255 60352 9271 60416
rect 9335 60352 9351 60416
rect 9415 60352 9423 60416
rect 9103 59328 9423 60352
rect 9103 59264 9111 59328
rect 9175 59264 9191 59328
rect 9255 59264 9271 59328
rect 9335 59264 9351 59328
rect 9415 59264 9423 59328
rect 9103 58240 9423 59264
rect 9103 58176 9111 58240
rect 9175 58176 9191 58240
rect 9255 58176 9271 58240
rect 9335 58176 9351 58240
rect 9415 58176 9423 58240
rect 9103 57152 9423 58176
rect 9103 57088 9111 57152
rect 9175 57088 9191 57152
rect 9255 57088 9271 57152
rect 9335 57088 9351 57152
rect 9415 57088 9423 57152
rect 9103 56064 9423 57088
rect 9103 56000 9111 56064
rect 9175 56000 9191 56064
rect 9255 56000 9271 56064
rect 9335 56000 9351 56064
rect 9415 56000 9423 56064
rect 9103 54976 9423 56000
rect 9103 54912 9111 54976
rect 9175 54912 9191 54976
rect 9255 54912 9271 54976
rect 9335 54912 9351 54976
rect 9415 54912 9423 54976
rect 9103 53888 9423 54912
rect 9103 53824 9111 53888
rect 9175 53824 9191 53888
rect 9255 53824 9271 53888
rect 9335 53824 9351 53888
rect 9415 53824 9423 53888
rect 9103 52800 9423 53824
rect 9103 52736 9111 52800
rect 9175 52736 9191 52800
rect 9255 52736 9271 52800
rect 9335 52736 9351 52800
rect 9415 52736 9423 52800
rect 9103 51712 9423 52736
rect 9103 51648 9111 51712
rect 9175 51648 9191 51712
rect 9255 51648 9271 51712
rect 9335 51648 9351 51712
rect 9415 51648 9423 51712
rect 9103 50624 9423 51648
rect 9103 50560 9111 50624
rect 9175 50560 9191 50624
rect 9255 50560 9271 50624
rect 9335 50560 9351 50624
rect 9415 50560 9423 50624
rect 9103 49536 9423 50560
rect 9103 49472 9111 49536
rect 9175 49472 9191 49536
rect 9255 49472 9271 49536
rect 9335 49472 9351 49536
rect 9415 49472 9423 49536
rect 9103 48448 9423 49472
rect 9103 48384 9111 48448
rect 9175 48384 9191 48448
rect 9255 48384 9271 48448
rect 9335 48384 9351 48448
rect 9415 48384 9423 48448
rect 9103 47360 9423 48384
rect 9103 47296 9111 47360
rect 9175 47296 9191 47360
rect 9255 47296 9271 47360
rect 9335 47296 9351 47360
rect 9415 47296 9423 47360
rect 9103 46272 9423 47296
rect 9103 46208 9111 46272
rect 9175 46208 9191 46272
rect 9255 46208 9271 46272
rect 9335 46208 9351 46272
rect 9415 46208 9423 46272
rect 9103 45184 9423 46208
rect 9103 45120 9111 45184
rect 9175 45120 9191 45184
rect 9255 45120 9271 45184
rect 9335 45120 9351 45184
rect 9415 45120 9423 45184
rect 9103 44096 9423 45120
rect 9103 44032 9111 44096
rect 9175 44032 9191 44096
rect 9255 44032 9271 44096
rect 9335 44032 9351 44096
rect 9415 44032 9423 44096
rect 9103 43008 9423 44032
rect 9103 42944 9111 43008
rect 9175 42944 9191 43008
rect 9255 42944 9271 43008
rect 9335 42944 9351 43008
rect 9415 42944 9423 43008
rect 9103 41920 9423 42944
rect 9103 41856 9111 41920
rect 9175 41856 9191 41920
rect 9255 41856 9271 41920
rect 9335 41856 9351 41920
rect 9415 41856 9423 41920
rect 9103 40832 9423 41856
rect 9103 40768 9111 40832
rect 9175 40768 9191 40832
rect 9255 40768 9271 40832
rect 9335 40768 9351 40832
rect 9415 40768 9423 40832
rect 9103 39744 9423 40768
rect 9103 39680 9111 39744
rect 9175 39680 9191 39744
rect 9255 39680 9271 39744
rect 9335 39680 9351 39744
rect 9415 39680 9423 39744
rect 9103 38656 9423 39680
rect 9103 38592 9111 38656
rect 9175 38592 9191 38656
rect 9255 38592 9271 38656
rect 9335 38592 9351 38656
rect 9415 38592 9423 38656
rect 9103 37568 9423 38592
rect 9103 37504 9111 37568
rect 9175 37504 9191 37568
rect 9255 37504 9271 37568
rect 9335 37504 9351 37568
rect 9415 37504 9423 37568
rect 9103 36480 9423 37504
rect 9103 36416 9111 36480
rect 9175 36416 9191 36480
rect 9255 36416 9271 36480
rect 9335 36416 9351 36480
rect 9415 36416 9423 36480
rect 9103 35392 9423 36416
rect 9103 35328 9111 35392
rect 9175 35328 9191 35392
rect 9255 35328 9271 35392
rect 9335 35328 9351 35392
rect 9415 35328 9423 35392
rect 9103 34304 9423 35328
rect 9103 34240 9111 34304
rect 9175 34240 9191 34304
rect 9255 34240 9271 34304
rect 9335 34240 9351 34304
rect 9415 34240 9423 34304
rect 9103 33216 9423 34240
rect 9103 33152 9111 33216
rect 9175 33152 9191 33216
rect 9255 33152 9271 33216
rect 9335 33152 9351 33216
rect 9415 33152 9423 33216
rect 9103 32128 9423 33152
rect 9103 32064 9111 32128
rect 9175 32064 9191 32128
rect 9255 32064 9271 32128
rect 9335 32064 9351 32128
rect 9415 32064 9423 32128
rect 9103 31040 9423 32064
rect 9103 30976 9111 31040
rect 9175 30976 9191 31040
rect 9255 30976 9271 31040
rect 9335 30976 9351 31040
rect 9415 30976 9423 31040
rect 9103 29952 9423 30976
rect 9103 29888 9111 29952
rect 9175 29888 9191 29952
rect 9255 29888 9271 29952
rect 9335 29888 9351 29952
rect 9415 29888 9423 29952
rect 9103 28864 9423 29888
rect 9103 28800 9111 28864
rect 9175 28800 9191 28864
rect 9255 28800 9271 28864
rect 9335 28800 9351 28864
rect 9415 28800 9423 28864
rect 9103 27776 9423 28800
rect 9103 27712 9111 27776
rect 9175 27712 9191 27776
rect 9255 27712 9271 27776
rect 9335 27712 9351 27776
rect 9415 27712 9423 27776
rect 9103 26688 9423 27712
rect 9103 26624 9111 26688
rect 9175 26624 9191 26688
rect 9255 26624 9271 26688
rect 9335 26624 9351 26688
rect 9415 26624 9423 26688
rect 9103 25600 9423 26624
rect 9103 25536 9111 25600
rect 9175 25536 9191 25600
rect 9255 25536 9271 25600
rect 9335 25536 9351 25600
rect 9415 25536 9423 25600
rect 9103 24512 9423 25536
rect 9103 24448 9111 24512
rect 9175 24448 9191 24512
rect 9255 24448 9271 24512
rect 9335 24448 9351 24512
rect 9415 24448 9423 24512
rect 9103 23424 9423 24448
rect 9103 23360 9111 23424
rect 9175 23360 9191 23424
rect 9255 23360 9271 23424
rect 9335 23360 9351 23424
rect 9415 23360 9423 23424
rect 9103 22336 9423 23360
rect 9103 22272 9111 22336
rect 9175 22272 9191 22336
rect 9255 22272 9271 22336
rect 9335 22272 9351 22336
rect 9415 22272 9423 22336
rect 9103 21248 9423 22272
rect 9103 21184 9111 21248
rect 9175 21184 9191 21248
rect 9255 21184 9271 21248
rect 9335 21184 9351 21248
rect 9415 21184 9423 21248
rect 9103 20160 9423 21184
rect 9103 20096 9111 20160
rect 9175 20096 9191 20160
rect 9255 20096 9271 20160
rect 9335 20096 9351 20160
rect 9415 20096 9423 20160
rect 9103 19072 9423 20096
rect 9103 19008 9111 19072
rect 9175 19008 9191 19072
rect 9255 19008 9271 19072
rect 9335 19008 9351 19072
rect 9415 19008 9423 19072
rect 9103 17984 9423 19008
rect 9103 17920 9111 17984
rect 9175 17920 9191 17984
rect 9255 17920 9271 17984
rect 9335 17920 9351 17984
rect 9415 17920 9423 17984
rect 9103 16896 9423 17920
rect 9103 16832 9111 16896
rect 9175 16832 9191 16896
rect 9255 16832 9271 16896
rect 9335 16832 9351 16896
rect 9415 16832 9423 16896
rect 9103 15808 9423 16832
rect 9103 15744 9111 15808
rect 9175 15744 9191 15808
rect 9255 15744 9271 15808
rect 9335 15744 9351 15808
rect 9415 15744 9423 15808
rect 9103 14720 9423 15744
rect 9103 14656 9111 14720
rect 9175 14656 9191 14720
rect 9255 14656 9271 14720
rect 9335 14656 9351 14720
rect 9415 14656 9423 14720
rect 9103 13632 9423 14656
rect 9103 13568 9111 13632
rect 9175 13568 9191 13632
rect 9255 13568 9271 13632
rect 9335 13568 9351 13632
rect 9415 13568 9423 13632
rect 9103 12544 9423 13568
rect 9103 12480 9111 12544
rect 9175 12480 9191 12544
rect 9255 12480 9271 12544
rect 9335 12480 9351 12544
rect 9415 12480 9423 12544
rect 9103 11456 9423 12480
rect 9103 11392 9111 11456
rect 9175 11392 9191 11456
rect 9255 11392 9271 11456
rect 9335 11392 9351 11456
rect 9415 11392 9423 11456
rect 9103 10368 9423 11392
rect 9103 10304 9111 10368
rect 9175 10304 9191 10368
rect 9255 10304 9271 10368
rect 9335 10304 9351 10368
rect 9415 10304 9423 10368
rect 9103 9280 9423 10304
rect 9103 9216 9111 9280
rect 9175 9216 9191 9280
rect 9255 9216 9271 9280
rect 9335 9216 9351 9280
rect 9415 9216 9423 9280
rect 9103 8192 9423 9216
rect 9103 8128 9111 8192
rect 9175 8128 9191 8192
rect 9255 8128 9271 8192
rect 9335 8128 9351 8192
rect 9415 8128 9423 8192
rect 9103 7104 9423 8128
rect 9103 7040 9111 7104
rect 9175 7040 9191 7104
rect 9255 7040 9271 7104
rect 9335 7040 9351 7104
rect 9415 7040 9423 7104
rect 9103 6016 9423 7040
rect 9103 5952 9111 6016
rect 9175 5952 9191 6016
rect 9255 5952 9271 6016
rect 9335 5952 9351 6016
rect 9415 5952 9423 6016
rect 9103 4928 9423 5952
rect 9103 4864 9111 4928
rect 9175 4864 9191 4928
rect 9255 4864 9271 4928
rect 9335 4864 9351 4928
rect 9415 4864 9423 4928
rect 9103 3840 9423 4864
rect 9103 3776 9111 3840
rect 9175 3776 9191 3840
rect 9255 3776 9271 3840
rect 9335 3776 9351 3840
rect 9415 3776 9423 3840
rect 9103 2752 9423 3776
rect 9103 2688 9111 2752
rect 9175 2688 9191 2752
rect 9255 2688 9271 2752
rect 9335 2688 9351 2752
rect 9415 2688 9423 2752
rect 9103 2128 9423 2688
use sky130_fd_sc_hd__decap_4  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635444444
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output122 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1635444444
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1635444444
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1635444444
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1635444444
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_19
timestamp 1635444444
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1635444444
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1635444444
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_31
timestamp 1635444444
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1635444444
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_43
timestamp 1635444444
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1635444444
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1635444444
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1635444444
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1635444444
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1635444444
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1635444444
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1635444444
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1635444444
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1635444444
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1635444444
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1635444444
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input120 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 10212 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input83
timestamp 1635444444
transform -1 0 10212 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1635444444
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1635444444
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635444444
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635444444
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1635444444
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635444444
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1635444444
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_14
timestamp 1635444444
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1635444444
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1635444444
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1635444444
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1635444444
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1635444444
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1635444444
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1635444444
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1635444444
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1635444444
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1635444444
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1635444444
transform 1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635444444
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1635444444
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635444444
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1635444444
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1635444444
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1635444444
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1635444444
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1635444444
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1635444444
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1635444444
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1635444444
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1635444444
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1635444444
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1635444444
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_93
timestamp 1635444444
transform 1 0 9660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1635444444
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1635444444
transform 1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635444444
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1635444444
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635444444
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1635444444
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_14
timestamp 1635444444
transform 1 0 2392 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1635444444
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _103_
timestamp 1635444444
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1635444444
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1635444444
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1635444444
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1635444444
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1635444444
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1635444444
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1635444444
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1635444444
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1635444444
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1635444444
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp 1635444444
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635444444
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1635444444
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635444444
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _097_
timestamp 1635444444
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1635444444
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_14
timestamp 1635444444
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_21
timestamp 1635444444
transform 1 0 3036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _099_
timestamp 1635444444
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_29
timestamp 1635444444
transform 1 0 3772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_34
timestamp 1635444444
transform 1 0 4232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 4232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_46
timestamp 1635444444
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1635444444
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1635444444
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1635444444
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1635444444
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1635444444
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_93
timestamp 1635444444
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1635444444
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1635444444
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635444444
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1635444444
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1635444444
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635444444
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635444444
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _095_
timestamp 1635444444
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _104_
timestamp 1635444444
transform -1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1635444444
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_14
timestamp 1635444444
transform 1 0 2392 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1635444444
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_13
timestamp 1635444444
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _094_
timestamp 1635444444
transform 1 0 2668 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkinv_2  _102_
timestamp 1635444444
transform -1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 1635444444
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1635444444
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1635444444
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_35
timestamp 1635444444
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1635444444
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _083_
timestamp 1635444444
transform -1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _096_
timestamp 1635444444
transform -1 0 4968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _100_
timestamp 1635444444
transform -1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1635444444
transform 1 0 4968 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1635444444
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1635444444
transform 1 0 6072 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1635444444
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1635444444
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1635444444
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1635444444
transform 1 0 7176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1635444444
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1635444444
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1635444444
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1635444444
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1635444444
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1635444444
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1635444444
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1635444444
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1635444444
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1635444444
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635444444
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635444444
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7
timestamp 1635444444
transform 1 0 1748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635444444
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1635444444
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1635444444
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _105_
timestamp 1635444444
transform -1 0 3220 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1635444444
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1635444444
transform 1 0 4048 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1635444444
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _110_
timestamp 1635444444
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1635444444
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1635444444
transform 1 0 6256 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1635444444
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1635444444
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1635444444
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1635444444
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1635444444
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1635444444
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1635444444
transform 1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635444444
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_11
timestamp 1635444444
transform 1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1635444444
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635444444
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 1635444444
transform 1 0 2852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _108_
timestamp 1635444444
transform 1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1635444444
transform -1 0 2852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_26
timestamp 1635444444
transform 1 0 3496 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_38
timestamp 1635444444
transform 1 0 4600 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1635444444
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1635444444
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1635444444
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1635444444
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1635444444
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1635444444
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1635444444
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635444444
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1635444444
transform 1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635444444
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _106_
timestamp 1635444444
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1635444444
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1635444444
transform 1 0 2392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1635444444
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _114_
timestamp 1635444444
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1635444444
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1635444444
transform 1 0 4048 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1635444444
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _120_
timestamp 1635444444
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1635444444
transform 1 0 5152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1635444444
transform 1 0 6256 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1635444444
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1635444444
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1635444444
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1635444444
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1635444444
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635444444
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1635444444
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635444444
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _112_
timestamp 1635444444
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1635444444
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_14
timestamp 1635444444
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_21
timestamp 1635444444
transform 1 0 3036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _118_
timestamp 1635444444
transform 1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _124_
timestamp 1635444444
transform 1 0 3404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_28
timestamp 1635444444
transform 1 0 3680 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_40
timestamp 1635444444
transform 1 0 4784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1635444444
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1635444444
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1635444444
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1635444444
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1635444444
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1635444444
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1635444444
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635444444
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_7
timestamp 1635444444
transform 1 0 1748 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635444444
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1635444444
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_16
timestamp 1635444444
transform 1 0 2576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1635444444
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _122_
timestamp 1635444444
transform -1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _126_
timestamp 1635444444
transform 1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1635444444
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1635444444
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1635444444
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1635444444
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1635444444
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1635444444
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1635444444
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1635444444
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1635444444
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1635444444
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 1635444444
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635444444
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_7
timestamp 1635444444
transform 1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_7
timestamp 1635444444
transform 1 0 1748 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635444444
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635444444
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1635444444
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1635444444
transform -1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1635444444
transform 1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1635444444
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_13
timestamp 1635444444
transform 1 0 2300 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1635444444
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _117_
timestamp 1635444444
transform -1 0 3312 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1635444444
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1635444444
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1635444444
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1635444444
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1635444444
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1635444444
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1635444444
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1635444444
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1635444444
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1635444444
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1635444444
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1635444444
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1635444444
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1635444444
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1635444444
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1635444444
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1635444444
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1635444444
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1635444444
transform 1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1635444444
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635444444
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635444444
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_7
timestamp 1635444444
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635444444
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1635444444
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_19
timestamp 1635444444
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_31
timestamp 1635444444
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_43
timestamp 1635444444
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1635444444
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1635444444
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1635444444
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1635444444
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1635444444
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_101
timestamp 1635444444
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_93
timestamp 1635444444
transform 1 0 9660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635444444
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_7
timestamp 1635444444
transform 1 0 1748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635444444
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1635444444
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1635444444
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1635444444
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1635444444
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1635444444
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1635444444
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1635444444
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1635444444
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1635444444
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1635444444
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1635444444
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1635444444
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1635444444
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635444444
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_7
timestamp 1635444444
transform 1 0 1748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635444444
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1635444444
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_19
timestamp 1635444444
transform 1 0 2852 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_31
timestamp 1635444444
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_43
timestamp 1635444444
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1635444444
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1635444444
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1635444444
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1635444444
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1635444444
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1635444444
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp 1635444444
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635444444
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_7
timestamp 1635444444
transform 1 0 1748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635444444
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1635444444
transform -1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1635444444
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1635444444
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1635444444
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1635444444
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1635444444
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1635444444
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1635444444
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1635444444
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1635444444
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1635444444
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1635444444
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_97
timestamp 1635444444
transform 1 0 10028 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635444444
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_7
timestamp 1635444444
transform 1 0 1748 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_7
timestamp 1635444444
transform 1 0 1748 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635444444
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635444444
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1635444444
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1635444444
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_15
timestamp 1635444444
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_13
timestamp 1635444444
transform 1 0 2300 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1635444444
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1635444444
transform 1 0 2392 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _150_
timestamp 1635444444
transform 1 0 2668 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1635444444
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1635444444
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1635444444
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1635444444
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1635444444
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1635444444
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1635444444
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1635444444
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1635444444
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1635444444
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1635444444
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1635444444
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1635444444
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1635444444
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1635444444
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1635444444
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1635444444
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1635444444
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_93
timestamp 1635444444
transform 1 0 9660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_97
timestamp 1635444444
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635444444
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635444444
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_7
timestamp 1635444444
transform 1 0 1748 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635444444
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1635444444
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1635444444
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _139_
timestamp 1635444444
transform -1 0 3588 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1635444444
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1635444444
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1635444444
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1635444444
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1635444444
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1635444444
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1635444444
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1635444444
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1635444444
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_93
timestamp 1635444444
transform 1 0 9660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635444444
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_7
timestamp 1635444444
transform 1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635444444
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _129_
timestamp 1635444444
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1635444444
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_14
timestamp 1635444444
transform 1 0 2392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1635444444
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _133_
timestamp 1635444444
transform 1 0 2760 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1635444444
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1635444444
transform 1 0 4048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1635444444
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _146_
timestamp 1635444444
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1635444444
transform 1 0 5152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1635444444
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1635444444
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1635444444
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1635444444
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1635444444
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp 1635444444
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635444444
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_7
timestamp 1635444444
transform 1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635444444
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _131_
timestamp 1635444444
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1635444444
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 1635444444
transform 1 0 2392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1635444444
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _137_
timestamp 1635444444
transform 1 0 2760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _144_
timestamp 1635444444
transform 1 0 3404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_28
timestamp 1635444444
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_40
timestamp 1635444444
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1635444444
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1635444444
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1635444444
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1635444444
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1635444444
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1635444444
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_93
timestamp 1635444444
transform 1 0 9660 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635444444
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_7
timestamp 1635444444
transform 1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635444444
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _135_
timestamp 1635444444
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1635444444
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_14
timestamp 1635444444
transform 1 0 2392 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1635444444
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _140_
timestamp 1635444444
transform 1 0 2760 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1635444444
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1635444444
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1635444444
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1635444444
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1635444444
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1635444444
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1635444444
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1635444444
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1635444444
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1635444444
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_97
timestamp 1635444444
transform 1 0 10028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635444444
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_7
timestamp 1635444444
transform 1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635444444
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _142_
timestamp 1635444444
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1635444444
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_14
timestamp 1635444444
transform 1 0 2392 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_21
timestamp 1635444444
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _148_
timestamp 1635444444
transform 1 0 2760 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_33
timestamp 1635444444
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1635444444
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1635444444
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1635444444
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1635444444
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1635444444
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1635444444
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1635444444
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_93
timestamp 1635444444
transform 1 0 9660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635444444
transform -1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_7
timestamp 1635444444
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_7
timestamp 1635444444
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635444444
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635444444
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _151_
timestamp 1635444444
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _155_
timestamp 1635444444
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1635444444
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1635444444
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_14
timestamp 1635444444
transform 1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1635444444
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_14
timestamp 1635444444
transform 1 0 2392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _153_
timestamp 1635444444
transform 1 0 2760 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1635444444
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1635444444
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_26
timestamp 1635444444
transform 1 0 3496 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_38
timestamp 1635444444
transform 1 0 4600 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1635444444
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1635444444
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1635444444
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1635444444
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1635444444
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1635444444
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1635444444
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1635444444
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1635444444
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1635444444
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1635444444
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1635444444
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1635444444
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_97
timestamp 1635444444
transform 1 0 10028 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_101
timestamp 1635444444
transform 1 0 10396 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_93
timestamp 1635444444
transform 1 0 9660 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635444444
transform -1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635444444
transform -1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_7
timestamp 1635444444
transform 1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635444444
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _157_
timestamp 1635444444
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1635444444
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_14
timestamp 1635444444
transform 1 0 2392 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1635444444
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1635444444
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1635444444
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1635444444
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1635444444
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1635444444
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1635444444
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1635444444
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1635444444
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1635444444
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1635444444
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635444444
transform -1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_7
timestamp 1635444444
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635444444
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _159_
timestamp 1635444444
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1635444444
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_14
timestamp 1635444444
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_26
timestamp 1635444444
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1635444444
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1635444444
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1635444444
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1635444444
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1635444444
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1635444444
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1635444444
transform 1 0 10396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_93
timestamp 1635444444
transform 1 0 9660 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635444444
transform -1 0 10856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_7
timestamp 1635444444
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635444444
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1635444444
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_19
timestamp 1635444444
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1635444444
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1635444444
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1635444444
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1635444444
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1635444444
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1635444444
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1635444444
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1635444444
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1635444444
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1635444444
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_97
timestamp 1635444444
transform 1 0 10028 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635444444
transform -1 0 10856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_7
timestamp 1635444444
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635444444
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1635444444
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_19
timestamp 1635444444
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_31
timestamp 1635444444
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_43
timestamp 1635444444
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1635444444
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1635444444
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1635444444
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1635444444
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1635444444
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_93
timestamp 1635444444
transform 1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 1635444444
transform 1 0 10212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1635444444
transform 1 0 9936 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635444444
transform -1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_7
timestamp 1635444444
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635444444
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1635444444
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1635444444
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1635444444
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1635444444
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1635444444
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1635444444
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1635444444
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1635444444
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1635444444
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1635444444
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1635444444
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1635444444
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1635444444
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1635444444
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1635444444
transform 1 0 9936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635444444
transform -1 0 10856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_7
timestamp 1635444444
transform 1 0 1748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_7
timestamp 1635444444
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635444444
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635444444
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1635444444
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1635444444
transform -1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_19
timestamp 1635444444
transform 1 0 2852 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1635444444
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_31
timestamp 1635444444
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1635444444
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1635444444
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1635444444
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_43
timestamp 1635444444
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1635444444
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1635444444
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1635444444
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1635444444
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1635444444
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1635444444
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1635444444
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1635444444
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1635444444
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1635444444
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp 1635444444
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_89
timestamp 1635444444
transform 1 0 9292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1635444444
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1635444444
transform -1 0 9292 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_93
timestamp 1635444444
transform 1 0 9660 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_99
timestamp 1635444444
transform 1 0 10212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1635444444
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9752 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9660 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635444444
transform -1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635444444
transform -1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_7
timestamp 1635444444
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635444444
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1635444444
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_19
timestamp 1635444444
transform 1 0 2852 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_25
timestamp 1635444444
transform 1 0 3404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _093_
timestamp 1635444444
transform -1 0 3404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_33
timestamp 1635444444
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1635444444
transform -1 0 4140 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1635444444
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1635444444
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1635444444
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1635444444
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1635444444
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_81
timestamp 1635444444
transform 1 0 8556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_88
timestamp 1635444444
transform 1 0 9200 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1635444444
transform -1 0 9200 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_99
timestamp 1635444444
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9568 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635444444
transform -1 0 10856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_11
timestamp 1635444444
transform 1 0 2116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1635444444
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635444444
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1635444444
transform -1 0 2116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_18
timestamp 1635444444
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _172_
timestamp 1635444444
transform 1 0 2484 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1635444444
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1635444444
transform 1 0 4048 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1635444444
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1635444444
transform 1 0 5152 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1635444444
transform 1 0 6256 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1635444444
transform 1 0 7360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1635444444
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1635444444
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_89
timestamp 1635444444
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1635444444
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1635444444
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 10212 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635444444
transform -1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_11
timestamp 1635444444
transform 1 0 2116 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1635444444
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635444444
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1635444444
transform -1 0 2116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _161_
timestamp 1635444444
transform 1 0 2668 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1635444444
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1635444444
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1635444444
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1635444444
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1635444444
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1635444444
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1635444444
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_81
timestamp 1635444444
transform 1 0 8556 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_87
timestamp 1635444444
transform 1 0 9108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1635444444
transform -1 0 9108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_99
timestamp 1635444444
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_2  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9476 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635444444
transform -1 0 10856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_11
timestamp 1635444444
transform 1 0 2116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1635444444
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635444444
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1635444444
transform -1 0 2116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_18
timestamp 1635444444
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _170_
timestamp 1635444444
transform 1 0 2484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1635444444
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1635444444
transform 1 0 4048 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1635444444
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _174_
timestamp 1635444444
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1635444444
transform 1 0 5152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1635444444
transform 1 0 6256 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1635444444
transform 1 0 7360 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1635444444
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1635444444
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1635444444
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1635444444
transform -1 0 9384 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_90
timestamp 1635444444
transform 1 0 9384 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_99
timestamp 1635444444
transform 1 0 10212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 10212 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635444444
transform -1 0 10856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_11
timestamp 1635444444
transform 1 0 2116 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1635444444
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1635444444
transform 1 0 2116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1635444444
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635444444
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635444444
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1635444444
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1635444444
transform -1 0 2116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_17
timestamp 1635444444
transform 1 0 2668 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_21
timestamp 1635444444
transform 1 0 3036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_18
timestamp 1635444444
transform 1 0 2760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _166_
timestamp 1635444444
transform 1 0 2484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _168_
timestamp 1635444444
transform 1 0 2760 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _176_
timestamp 1635444444
transform 1 0 3404 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_28
timestamp 1635444444
transform 1 0 3680 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1635444444
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1635444444
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1635444444
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_40
timestamp 1635444444
transform 1 0 4784 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1635444444
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1635444444
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1635444444
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1635444444
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1635444444
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1635444444
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1635444444
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1635444444
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1635444444
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1635444444
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1635444444
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1635444444
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_93
timestamp 1635444444
transform 1 0 9660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_99
timestamp 1635444444
transform 1 0 10212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1635444444
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1635444444
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _084_
timestamp 1635444444
transform 1 0 9936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1635444444
transform 1 0 9936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635444444
transform -1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635444444
transform -1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_11
timestamp 1635444444
transform 1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1635444444
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635444444
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1635444444
transform -1 0 2116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_18
timestamp 1635444444
transform 1 0 2760 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_25
timestamp 1635444444
transform 1 0 3404 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _162_
timestamp 1635444444
transform 1 0 2484 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _164_
timestamp 1635444444
transform 1 0 3128 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_37
timestamp 1635444444
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1635444444
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1635444444
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1635444444
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1635444444
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1635444444
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1635444444
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_93
timestamp 1635444444
transform 1 0 9660 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1635444444
transform 1 0 10212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1635444444
transform 1 0 9936 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635444444
transform -1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_11
timestamp 1635444444
transform 1 0 2116 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1635444444
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635444444
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1635444444
transform -1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_23
timestamp 1635444444
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1635444444
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1635444444
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1635444444
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1635444444
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1635444444
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1635444444
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1635444444
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1635444444
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1635444444
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1635444444
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_93
timestamp 1635444444
transform 1 0 9660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1635444444
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1635444444
transform 1 0 9936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635444444
transform -1 0 10856 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_11
timestamp 1635444444
transform 1 0 2116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1635444444
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635444444
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1635444444
transform -1 0 2116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_23
timestamp 1635444444
transform 1 0 3220 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_35
timestamp 1635444444
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1635444444
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1635444444
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1635444444
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1635444444
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1635444444
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1635444444
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_93
timestamp 1635444444
transform 1 0 9660 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_99
timestamp 1635444444
transform 1 0 10212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _088_
timestamp 1635444444
transform 1 0 9752 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635444444
transform -1 0 10856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_11
timestamp 1635444444
transform 1 0 2116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1635444444
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635444444
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1635444444
transform -1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_23
timestamp 1635444444
transform 1 0 3220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1635444444
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1635444444
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1635444444
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1635444444
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1635444444
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1635444444
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1635444444
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1635444444
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_85
timestamp 1635444444
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1635444444
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_99
timestamp 1635444444
transform 1 0 10212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _090_
timestamp 1635444444
transform -1 0 10212 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635444444
transform -1 0 10856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1635444444
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635444444
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1635444444
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1635444444
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1635444444
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1635444444
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1635444444
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1635444444
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1635444444
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1635444444
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1635444444
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_93
timestamp 1635444444
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_99
timestamp 1635444444
transform 1 0 10212 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1635444444
transform 1 0 9936 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635444444
transform -1 0 10856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_11
timestamp 1635444444
transform 1 0 2116 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1635444444
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_7
timestamp 1635444444
transform 1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635444444
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1635444444
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _183_
timestamp 1635444444
transform 1 0 2116 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1635444444
transform -1 0 2116 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input33
timestamp 1635444444
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 1635444444
transform 1 0 3220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_14
timestamp 1635444444
transform 1 0 2392 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_21
timestamp 1635444444
transform 1 0 3036 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _185_
timestamp 1635444444
transform 1 0 2760 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1635444444
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1635444444
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_33
timestamp 1635444444
transform 1 0 4140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1635444444
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1635444444
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_45
timestamp 1635444444
transform 1 0 5244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1635444444
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1635444444
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1635444444
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1635444444
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1635444444
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1635444444
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1635444444
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1635444444
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1635444444
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1635444444
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1635444444
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_93
timestamp 1635444444
transform 1 0 9660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1635444444
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_93
timestamp 1635444444
transform 1 0 9660 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_99
timestamp 1635444444
transform 1 0 10212 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1635444444
transform 1 0 9936 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1635444444
transform 1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635444444
transform -1 0 10856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1635444444
transform -1 0 10856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_7
timestamp 1635444444
transform 1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1635444444
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _181_
timestamp 1635444444
transform 1 0 2116 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1635444444
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_14
timestamp 1635444444
transform 1 0 2392 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1635444444
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _182_
timestamp 1635444444
transform 1 0 2760 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1635444444
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1635444444
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1635444444
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1635444444
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1635444444
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1635444444
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1635444444
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1635444444
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1635444444
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1635444444
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_93
timestamp 1635444444
transform 1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_99
timestamp 1635444444
transform 1 0 10212 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1635444444
transform 1 0 9936 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1635444444
transform -1 0 10856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_7
timestamp 1635444444
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1635444444
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _184_
timestamp 1635444444
transform 1 0 2116 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1635444444
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_14
timestamp 1635444444
transform 1 0 2392 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_26
timestamp 1635444444
transform 1 0 3496 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_38
timestamp 1635444444
transform 1 0 4600 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_50
timestamp 1635444444
transform 1 0 5704 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1635444444
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1635444444
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1635444444
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1635444444
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_89
timestamp 1635444444
transform 1 0 9292 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_99
timestamp 1635444444
transform 1 0 10212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_1  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9384 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1635444444
transform -1 0 10856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_7
timestamp 1635444444
transform 1 0 1748 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1635444444
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1635444444
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1635444444
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _186_
timestamp 1635444444
transform 1 0 2300 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1635444444
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1635444444
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1635444444
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1635444444
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1635444444
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1635444444
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1635444444
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1635444444
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1635444444
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1635444444
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_93
timestamp 1635444444
transform 1 0 9660 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_99
timestamp 1635444444
transform 1 0 10212 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1635444444
transform 1 0 9936 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1635444444
transform -1 0 10856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_7
timestamp 1635444444
transform 1 0 1748 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1635444444
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1635444444
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_15
timestamp 1635444444
transform 1 0 2484 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _180_
timestamp 1635444444
transform 1 0 2576 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_51_26
timestamp 1635444444
transform 1 0 3496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_34
timestamp 1635444444
transform 1 0 4232 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _107_
timestamp 1635444444
transform -1 0 4232 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_46
timestamp 1635444444
transform 1 0 5336 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1635444444
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1635444444
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1635444444
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1635444444
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1635444444
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_93
timestamp 1635444444
transform 1 0 9660 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_99
timestamp 1635444444
transform 1 0 10212 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1635444444
transform 1 0 9936 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1635444444
transform -1 0 10856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_7
timestamp 1635444444
transform 1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_7
timestamp 1635444444
transform 1 0 1748 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1635444444
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1635444444
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _187_
timestamp 1635444444
transform 1 0 2116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _188_
timestamp 1635444444
transform 1 0 2116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1635444444
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1635444444
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_14
timestamp 1635444444
transform 1 0 2392 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1635444444
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_14
timestamp 1635444444
transform 1 0 2392 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_20
timestamp 1635444444
transform 1 0 2944 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_25
timestamp 1635444444
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _111_
timestamp 1635444444
transform -1 0 3404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _189_
timestamp 1635444444
transform 1 0 2760 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1635444444
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_33
timestamp 1635444444
transform 1 0 4140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_37
timestamp 1635444444
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1635444444
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _109_
timestamp 1635444444
transform -1 0 4140 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_45
timestamp 1635444444
transform 1 0 5244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_49
timestamp 1635444444
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_57
timestamp 1635444444
transform 1 0 6348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1635444444
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1635444444
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1635444444
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_69
timestamp 1635444444
transform 1 0 7452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1635444444
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_81
timestamp 1635444444
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1635444444
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1635444444
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1635444444
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_93
timestamp 1635444444
transform 1 0 9660 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1635444444
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_93
timestamp 1635444444
transform 1 0 9660 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_99
timestamp 1635444444
transform 1 0 10212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1635444444
transform 1 0 9936 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1635444444
transform 1 0 9936 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1635444444
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1635444444
transform -1 0 10856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_7
timestamp 1635444444
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1635444444
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _190_
timestamp 1635444444
transform 1 0 2116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1635444444
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_14
timestamp 1635444444
transform 1 0 2392 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1635444444
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _113_
timestamp 1635444444
transform -1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1635444444
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1635444444
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1635444444
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1635444444
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1635444444
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1635444444
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1635444444
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1635444444
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1635444444
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_97
timestamp 1635444444
transform 1 0 10028 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1635444444
transform -1 0 10856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_7
timestamp 1635444444
transform 1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1635444444
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _191_
timestamp 1635444444
transform 1 0 2116 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1635444444
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_14
timestamp 1635444444
transform 1 0 2392 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_26
timestamp 1635444444
transform 1 0 3496 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_38
timestamp 1635444444
transform 1 0 4600 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_50
timestamp 1635444444
transform 1 0 5704 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1635444444
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1635444444
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1635444444
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1635444444
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_93
timestamp 1635444444
transform 1 0 9660 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_99
timestamp 1635444444
transform 1 0 10212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1635444444
transform 1 0 9936 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1635444444
transform -1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_7
timestamp 1635444444
transform 1 0 1748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1635444444
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1635444444
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_19
timestamp 1635444444
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1635444444
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1635444444
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1635444444
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1635444444
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1635444444
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1635444444
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1635444444
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1635444444
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1635444444
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1635444444
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_93
timestamp 1635444444
transform 1 0 9660 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_99
timestamp 1635444444
transform 1 0 10212 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1635444444
transform 1 0 9936 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1635444444
transform -1 0 10856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_7
timestamp 1635444444
transform 1 0 1748 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1635444444
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1635444444
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_19
timestamp 1635444444
transform 1 0 2852 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_31
timestamp 1635444444
transform 1 0 3956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_43
timestamp 1635444444
transform 1 0 5060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1635444444
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1635444444
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1635444444
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1635444444
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1635444444
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_101
timestamp 1635444444
transform 1 0 10396 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_93
timestamp 1635444444
transform 1 0 9660 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1635444444
transform -1 0 10856 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_7
timestamp 1635444444
transform 1 0 1748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1635444444
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1635444444
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 1635444444
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1635444444
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1635444444
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1635444444
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1635444444
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1635444444
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1635444444
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1635444444
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1635444444
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1635444444
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1635444444
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_93
timestamp 1635444444
transform 1 0 9660 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_99
timestamp 1635444444
transform 1 0 10212 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1635444444
transform 1 0 9936 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1635444444
transform -1 0 10856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_7
timestamp 1635444444
transform 1 0 1748 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_7
timestamp 1635444444
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1635444444
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1635444444
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1635444444
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1635444444
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_19
timestamp 1635444444
transform 1 0 2852 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 1635444444
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_31
timestamp 1635444444
transform 1 0 3956 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_36
timestamp 1635444444
transform 1 0 4416 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1635444444
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_29
timestamp 1635444444
transform 1 0 3772 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_36
timestamp 1635444444
transform 1 0 4416 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1635444444
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _115_
timestamp 1635444444
transform -1 0 4416 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _119_
timestamp 1635444444
transform -1 0 4416 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_48
timestamp 1635444444
transform 1 0 5520 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_48
timestamp 1635444444
transform 1 0 5520 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1635444444
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_60
timestamp 1635444444
transform 1 0 6624 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1635444444
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1635444444
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_72
timestamp 1635444444
transform 1 0 7728 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1635444444
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_85
timestamp 1635444444
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1635444444
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_93
timestamp 1635444444
transform 1 0 9660 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_99
timestamp 1635444444
transform 1 0 10212 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_93
timestamp 1635444444
transform 1 0 9660 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_99
timestamp 1635444444
transform 1 0 10212 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1635444444
transform 1 0 9936 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1635444444
transform 1 0 9936 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1635444444
transform -1 0 10856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1635444444
transform -1 0 10856 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1635444444
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1635444444
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _196_
timestamp 1635444444
transform 1 0 2116 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1635444444
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_14
timestamp 1635444444
transform 1 0 2392 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_26
timestamp 1635444444
transform 1 0 3496 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_36
timestamp 1635444444
transform 1 0 4416 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _121_
timestamp 1635444444
transform -1 0 4416 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_48
timestamp 1635444444
transform 1 0 5520 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1635444444
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1635444444
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1635444444
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1635444444
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_101
timestamp 1635444444
transform 1 0 10396 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_93
timestamp 1635444444
transform 1 0 9660 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1635444444
transform -1 0 10856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_7
timestamp 1635444444
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1635444444
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _194_
timestamp 1635444444
transform 1 0 2116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1635444444
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_14
timestamp 1635444444
transform 1 0 2392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1635444444
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _195_
timestamp 1635444444
transform 1 0 2760 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1635444444
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_29
timestamp 1635444444
transform 1 0 3772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_36
timestamp 1635444444
transform 1 0 4416 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1635444444
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _123_
timestamp 1635444444
transform -1 0 4416 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_48
timestamp 1635444444
transform 1 0 5520 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_60
timestamp 1635444444
transform 1 0 6624 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_72
timestamp 1635444444
transform 1 0 7728 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_85
timestamp 1635444444
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1635444444
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_93
timestamp 1635444444
transform 1 0 9660 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_99
timestamp 1635444444
transform 1 0 10212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1635444444
transform 1 0 9936 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1635444444
transform -1 0 10856 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_7
timestamp 1635444444
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1635444444
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _197_
timestamp 1635444444
transform 1 0 2116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1635444444
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_14
timestamp 1635444444
transform 1 0 2392 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_21
timestamp 1635444444
transform 1 0 3036 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _198_
timestamp 1635444444
transform 1 0 2760 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_29
timestamp 1635444444
transform 1 0 3772 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_36
timestamp 1635444444
transform 1 0 4416 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _125_
timestamp 1635444444
transform -1 0 4416 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_48
timestamp 1635444444
transform 1 0 5520 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1635444444
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1635444444
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1635444444
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1635444444
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_93
timestamp 1635444444
transform 1 0 9660 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_99
timestamp 1635444444
transform 1 0 10212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1635444444
transform 1 0 9936 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1635444444
transform -1 0 10856 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_7
timestamp 1635444444
transform 1 0 1748 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1635444444
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1635444444
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_13
timestamp 1635444444
transform 1 0 2300 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1635444444
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _193_
timestamp 1635444444
transform 1 0 2392 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_64_33
timestamp 1635444444
transform 1 0 4140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1635444444
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _127_
timestamp 1635444444
transform -1 0 4140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_45
timestamp 1635444444
transform 1 0 5244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_57
timestamp 1635444444
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_69
timestamp 1635444444
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1635444444
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1635444444
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1635444444
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_93
timestamp 1635444444
transform 1 0 9660 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_99
timestamp 1635444444
transform 1 0 10212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1635444444
transform 1 0 9936 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1635444444
transform -1 0 10856 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_7
timestamp 1635444444
transform 1 0 1748 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1635444444
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1635444444
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_13
timestamp 1635444444
transform 1 0 2300 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_24
timestamp 1635444444
transform 1 0 3312 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _199_
timestamp 1635444444
transform 1 0 2392 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_65_32
timestamp 1635444444
transform 1 0 4048 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _130_
timestamp 1635444444
transform -1 0 4048 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_44
timestamp 1635444444
transform 1 0 5152 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1635444444
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1635444444
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1635444444
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1635444444
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_101
timestamp 1635444444
transform 1 0 10396 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_93
timestamp 1635444444
transform 1 0 9660 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1635444444
transform -1 0 10856 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_7
timestamp 1635444444
transform 1 0 1748 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_7
timestamp 1635444444
transform 1 0 1748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1635444444
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1635444444
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _200_
timestamp 1635444444
transform 1 0 2116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _201_
timestamp 1635444444
transform 1 0 2116 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1635444444
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1635444444
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_14
timestamp 1635444444
transform 1 0 2392 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_21
timestamp 1635444444
transform 1 0 3036 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_14
timestamp 1635444444
transform 1 0 2392 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_21
timestamp 1635444444
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _202_
timestamp 1635444444
transform 1 0 2760 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _204_
timestamp 1635444444
transform 1 0 2760 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1635444444
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_33
timestamp 1635444444
transform 1 0 4140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_33
timestamp 1635444444
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1635444444
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _132_
timestamp 1635444444
transform -1 0 4140 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_45
timestamp 1635444444
transform 1 0 5244 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1635444444
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_57
timestamp 1635444444
transform 1 0 6348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1635444444
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1635444444
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1635444444
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_69
timestamp 1635444444
transform 1 0 7452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1635444444
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_81
timestamp 1635444444
transform 1 0 8556 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_85
timestamp 1635444444
transform 1 0 8924 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1635444444
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1635444444
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_93
timestamp 1635444444
transform 1 0 9660 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_99
timestamp 1635444444
transform 1 0 10212 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_93
timestamp 1635444444
transform 1 0 9660 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_99
timestamp 1635444444
transform 1 0 10212 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1635444444
transform 1 0 9936 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1635444444
transform 1 0 9936 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1635444444
transform -1 0 10856 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1635444444
transform -1 0 10856 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_7
timestamp 1635444444
transform 1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1635444444
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _203_
timestamp 1635444444
transform 1 0 2116 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1635444444
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_14
timestamp 1635444444
transform 1 0 2392 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_26
timestamp 1635444444
transform 1 0 3496 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_33
timestamp 1635444444
transform 1 0 4140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1635444444
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _134_
timestamp 1635444444
transform -1 0 4140 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_45
timestamp 1635444444
transform 1 0 5244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_57
timestamp 1635444444
transform 1 0 6348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_69
timestamp 1635444444
transform 1 0 7452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_81
timestamp 1635444444
transform 1 0 8556 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1635444444
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1635444444
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_97
timestamp 1635444444
transform 1 0 10028 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1635444444
transform -1 0 10856 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_7
timestamp 1635444444
transform 1 0 1748 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1635444444
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1635444444
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_15
timestamp 1635444444
transform 1 0 2484 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _205_
timestamp 1635444444
transform 1 0 2576 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_69_26
timestamp 1635444444
transform 1 0 3496 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_34
timestamp 1635444444
transform 1 0 4232 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _136_
timestamp 1635444444
transform -1 0 4232 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_46
timestamp 1635444444
transform 1 0 5336 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_54
timestamp 1635444444
transform 1 0 6072 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1635444444
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1635444444
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1635444444
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1635444444
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_93
timestamp 1635444444
transform 1 0 9660 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_99
timestamp 1635444444
transform 1 0 10212 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1635444444
transform 1 0 9936 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1635444444
transform -1 0 10856 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_7
timestamp 1635444444
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1635444444
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _206_
timestamp 1635444444
transform 1 0 2116 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1635444444
transform -1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_14
timestamp 1635444444
transform 1 0 2392 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_21
timestamp 1635444444
transform 1 0 3036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 1635444444
transform 1 0 2760 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1635444444
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_29
timestamp 1635444444
transform 1 0 3772 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_34
timestamp 1635444444
transform 1 0 4232 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1635444444
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _138_
timestamp 1635444444
transform -1 0 4232 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_46
timestamp 1635444444
transform 1 0 5336 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_58
timestamp 1635444444
transform 1 0 6440 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_70
timestamp 1635444444
transform 1 0 7544 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_82
timestamp 1635444444
transform 1 0 8648 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_85
timestamp 1635444444
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1635444444
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_93
timestamp 1635444444
transform 1 0 9660 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_99
timestamp 1635444444
transform 1 0 10212 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1635444444
transform 1 0 9936 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1635444444
transform -1 0 10856 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_7
timestamp 1635444444
transform 1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1635444444
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _208_
timestamp 1635444444
transform 1 0 2116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1635444444
transform -1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_14
timestamp 1635444444
transform 1 0 2392 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_21
timestamp 1635444444
transform 1 0 3036 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _209_
timestamp 1635444444
transform 1 0 2760 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_71_29
timestamp 1635444444
transform 1 0 3772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_34
timestamp 1635444444
transform 1 0 4232 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _141_
timestamp 1635444444
transform -1 0 4232 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_46
timestamp 1635444444
transform 1 0 5336 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp 1635444444
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1635444444
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1635444444
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1635444444
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1635444444
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_93
timestamp 1635444444
transform 1 0 9660 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_99
timestamp 1635444444
transform 1 0 10212 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1635444444
transform 1 0 9936 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1635444444
transform -1 0 10856 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_7
timestamp 1635444444
transform 1 0 1748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_7
timestamp 1635444444
transform 1 0 1748 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1635444444
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1635444444
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _210_
timestamp 1635444444
transform 1 0 2116 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1635444444
transform -1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1635444444
transform -1 0 1748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_14
timestamp 1635444444
transform 1 0 2392 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_19
timestamp 1635444444
transform 1 0 2852 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_26
timestamp 1635444444
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_33
timestamp 1635444444
transform 1 0 4140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_27
timestamp 1635444444
transform 1 0 3588 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_32
timestamp 1635444444
transform 1 0 4048 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1635444444
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _143_
timestamp 1635444444
transform -1 0 4140 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _145_
timestamp 1635444444
transform -1 0 4048 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_45
timestamp 1635444444
transform 1 0 5244 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_44
timestamp 1635444444
transform 1 0 5152 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_57
timestamp 1635444444
transform 1 0 6348 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1635444444
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1635444444
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_69
timestamp 1635444444
transform 1 0 7452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1635444444
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_81
timestamp 1635444444
transform 1 0 8556 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1635444444
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1635444444
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1635444444
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_97
timestamp 1635444444
transform 1 0 10028 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_73_93
timestamp 1635444444
transform 1 0 9660 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_99
timestamp 1635444444
transform 1 0 10212 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1635444444
transform 1 0 9936 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1635444444
transform -1 0 10856 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1635444444
transform -1 0 10856 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_7
timestamp 1635444444
transform 1 0 1748 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1635444444
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1635444444
transform -1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_19
timestamp 1635444444
transform 1 0 2852 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1635444444
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1635444444
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _192_
timestamp 1635444444
transform 1 0 3772 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_74_39
timestamp 1635444444
transform 1 0 4692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_51
timestamp 1635444444
transform 1 0 5796 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_63
timestamp 1635444444
transform 1 0 6900 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_75
timestamp 1635444444
transform 1 0 8004 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1635444444
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_85
timestamp 1635444444
transform 1 0 8924 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1635444444
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_93
timestamp 1635444444
transform 1 0 9660 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_99
timestamp 1635444444
transform 1 0 10212 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1635444444
transform 1 0 9936 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1635444444
transform -1 0 10856 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_7
timestamp 1635444444
transform 1 0 1748 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1635444444
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1635444444
transform -1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_19
timestamp 1635444444
transform 1 0 2852 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_25
timestamp 1635444444
transform 1 0 3404 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_30
timestamp 1635444444
transform 1 0 3864 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _147_
timestamp 1635444444
transform -1 0 3864 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_42
timestamp 1635444444
transform 1 0 4968 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_54
timestamp 1635444444
transform 1 0 6072 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1635444444
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1635444444
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1635444444
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1635444444
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_101
timestamp 1635444444
transform 1 0 10396 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_93
timestamp 1635444444
transform 1 0 9660 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1635444444
transform -1 0 10856 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_7
timestamp 1635444444
transform 1 0 1748 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1635444444
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1635444444
transform -1 0 1748 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_19
timestamp 1635444444
transform 1 0 2852 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1635444444
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1635444444
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1635444444
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1635444444
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1635444444
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1635444444
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1635444444
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1635444444
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_85
timestamp 1635444444
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1635444444
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_93
timestamp 1635444444
transform 1 0 9660 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_99
timestamp 1635444444
transform 1 0 10212 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1635444444
transform 1 0 9936 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1635444444
transform -1 0 10856 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_7
timestamp 1635444444
transform 1 0 1748 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1635444444
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1635444444
transform -1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_19
timestamp 1635444444
transform 1 0 2852 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_31
timestamp 1635444444
transform 1 0 3956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_43
timestamp 1635444444
transform 1 0 5060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1635444444
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1635444444
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1635444444
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1635444444
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1635444444
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_93
timestamp 1635444444
transform 1 0 9660 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_99
timestamp 1635444444
transform 1 0 10212 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1635444444
transform 1 0 9936 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1635444444
transform -1 0 10856 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_7
timestamp 1635444444
transform 1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1635444444
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _212_
timestamp 1635444444
transform 1 0 2116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1635444444
transform -1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_14
timestamp 1635444444
transform 1 0 2392 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_21
timestamp 1635444444
transform 1 0 3036 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _214_
timestamp 1635444444
transform 1 0 2760 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1635444444
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_29
timestamp 1635444444
transform 1 0 3772 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_35
timestamp 1635444444
transform 1 0 4324 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1635444444
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _149_
timestamp 1635444444
transform -1 0 4324 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_47
timestamp 1635444444
transform 1 0 5428 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_59
timestamp 1635444444
transform 1 0 6532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_71
timestamp 1635444444
transform 1 0 7636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1635444444
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_85
timestamp 1635444444
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1635444444
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_93
timestamp 1635444444
transform 1 0 9660 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_99
timestamp 1635444444
transform 1 0 10212 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1635444444
transform 1 0 9936 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1635444444
transform -1 0 10856 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_7
timestamp 1635444444
transform 1 0 1748 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_7
timestamp 1635444444
transform 1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1635444444
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1635444444
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _213_
timestamp 1635444444
transform 1 0 2116 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1635444444
transform -1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1635444444
transform -1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_15
timestamp 1635444444
transform 1 0 2484 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_14
timestamp 1635444444
transform 1 0 2392 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1635444444
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _211_
timestamp 1635444444
transform 1 0 2668 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _215_
timestamp 1635444444
transform -1 0 3036 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_27
timestamp 1635444444
transform 1 0 3588 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_35
timestamp 1635444444
transform 1 0 4324 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1635444444
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_33
timestamp 1635444444
transform 1 0 4140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1635444444
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _152_
timestamp 1635444444
transform -1 0 4324 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _154_
timestamp 1635444444
transform -1 0 4140 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_47
timestamp 1635444444
transform 1 0 5428 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_45
timestamp 1635444444
transform 1 0 5244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1635444444
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1635444444
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_57
timestamp 1635444444
transform 1 0 6348 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1635444444
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1635444444
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_69
timestamp 1635444444
transform 1 0 7452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1635444444
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_81
timestamp 1635444444
transform 1 0 8556 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_85
timestamp 1635444444
transform 1 0 8924 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1635444444
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_101
timestamp 1635444444
transform 1 0 10396 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_93
timestamp 1635444444
transform 1 0 9660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_93
timestamp 1635444444
transform 1 0 9660 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_99
timestamp 1635444444
transform 1 0 10212 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1635444444
transform 1 0 9936 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1635444444
transform -1 0 10856 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1635444444
transform -1 0 10856 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_7
timestamp 1635444444
transform 1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1635444444
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _216_
timestamp 1635444444
transform 1 0 2116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1635444444
transform -1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_14
timestamp 1635444444
transform 1 0 2392 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_22
timestamp 1635444444
transform 1 0 3128 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _156_
timestamp 1635444444
transform -1 0 3772 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_29
timestamp 1635444444
transform 1 0 3772 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_41
timestamp 1635444444
transform 1 0 4876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_53
timestamp 1635444444
transform 1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1635444444
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1635444444
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1635444444
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1635444444
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_93
timestamp 1635444444
transform 1 0 9660 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_99
timestamp 1635444444
transform 1 0 10212 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1635444444
transform 1 0 9936 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1635444444
transform -1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_7
timestamp 1635444444
transform 1 0 1748 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1635444444
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1635444444
transform -1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_19
timestamp 1635444444
transform 1 0 2852 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1635444444
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1635444444
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1635444444
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1635444444
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1635444444
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1635444444
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1635444444
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1635444444
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_85
timestamp 1635444444
transform 1 0 8924 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1635444444
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_93
timestamp 1635444444
transform 1 0 9660 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_99
timestamp 1635444444
transform 1 0 10212 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1635444444
transform 1 0 9936 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1635444444
transform -1 0 10856 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_7
timestamp 1635444444
transform 1 0 1748 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1635444444
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1635444444
transform -1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_83_15
timestamp 1635444444
transform 1 0 2484 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _217_
timestamp 1635444444
transform -1 0 3680 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_83_28
timestamp 1635444444
transform 1 0 3680 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_36
timestamp 1635444444
transform 1 0 4416 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _158_
timestamp 1635444444
transform -1 0 4416 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_48
timestamp 1635444444
transform 1 0 5520 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1635444444
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1635444444
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1635444444
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1635444444
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_101
timestamp 1635444444
transform 1 0 10396 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_93
timestamp 1635444444
transform 1 0 9660 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1635444444
transform -1 0 10856 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_7
timestamp 1635444444
transform 1 0 1748 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1635444444
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1635444444
transform -1 0 1748 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_19
timestamp 1635444444
transform 1 0 2852 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1635444444
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1635444444
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1635444444
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1635444444
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1635444444
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1635444444
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1635444444
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1635444444
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_85
timestamp 1635444444
transform 1 0 8924 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1635444444
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_84_93
timestamp 1635444444
transform 1 0 9660 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_99
timestamp 1635444444
transform 1 0 10212 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1635444444
transform 1 0 9936 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1635444444
transform -1 0 10856 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_7
timestamp 1635444444
transform 1 0 1748 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_7
timestamp 1635444444
transform 1 0 1748 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1635444444
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1635444444
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1635444444
transform -1 0 1748 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1635444444
transform -1 0 1748 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_19
timestamp 1635444444
transform 1 0 2852 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_16
timestamp 1635444444
transform 1 0 2576 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _218_
timestamp 1635444444
transform 1 0 2300 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_85_27
timestamp 1635444444
transform 1 0 3588 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_32
timestamp 1635444444
transform 1 0 4048 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_29
timestamp 1635444444
transform 1 0 3772 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_35
timestamp 1635444444
transform 1 0 4324 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1635444444
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _160_
timestamp 1635444444
transform -1 0 4324 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _229_
timestamp 1635444444
transform -1 0 4048 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_44
timestamp 1635444444
transform 1 0 5152 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_47
timestamp 1635444444
transform 1 0 5428 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1635444444
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_59
timestamp 1635444444
transform 1 0 6532 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1635444444
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1635444444
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_71
timestamp 1635444444
transform 1 0 7636 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1635444444
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1635444444
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_85
timestamp 1635444444
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1635444444
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_93
timestamp 1635444444
transform 1 0 9660 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_99
timestamp 1635444444
transform 1 0 10212 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_97
timestamp 1635444444
transform 1 0 10028 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1635444444
transform 1 0 9936 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1635444444
transform -1 0 10856 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1635444444
transform -1 0 10856 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_87_7
timestamp 1635444444
transform 1 0 1748 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1635444444
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1635444444
transform -1 0 1748 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_16
timestamp 1635444444
transform 1 0 2576 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _179_
timestamp 1635444444
transform -1 0 3496 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _219_
timestamp 1635444444
transform 1 0 2300 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_26
timestamp 1635444444
transform 1 0 3496 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_30
timestamp 1635444444
transform 1 0 3864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_35
timestamp 1635444444
transform 1 0 4324 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _163_
timestamp 1635444444
transform -1 0 4324 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_47
timestamp 1635444444
transform 1 0 5428 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1635444444
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1635444444
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1635444444
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1635444444
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1635444444
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_93
timestamp 1635444444
transform 1 0 9660 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_99
timestamp 1635444444
transform 1 0 10212 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1635444444
transform 1 0 9936 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1635444444
transform -1 0 10856 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_10
timestamp 1635444444
transform 1 0 2024 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1635444444
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_88_18
timestamp 1635444444
transform 1 0 2760 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1635444444
transform -1 0 2760 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1635444444
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_29
timestamp 1635444444
transform 1 0 3772 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_88_35
timestamp 1635444444
transform 1 0 4324 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1635444444
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _165_
timestamp 1635444444
transform -1 0 4324 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_47
timestamp 1635444444
transform 1 0 5428 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_59
timestamp 1635444444
transform 1 0 6532 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_71
timestamp 1635444444
transform 1 0 7636 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1635444444
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_85
timestamp 1635444444
transform 1 0 8924 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1635444444
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_93
timestamp 1635444444
transform 1 0 9660 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_99
timestamp 1635444444
transform 1 0 10212 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1635444444
transform 1 0 9936 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1635444444
transform -1 0 10856 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_10
timestamp 1635444444
transform 1 0 2024 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1635444444
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _234_
timestamp 1635444444
transform 1 0 1380 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_89_18
timestamp 1635444444
transform 1 0 2760 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_25
timestamp 1635444444
transform 1 0 3404 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _220_
timestamp 1635444444
transform 1 0 3128 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1635444444
transform 1 0 2392 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_35
timestamp 1635444444
transform 1 0 4324 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _167_
timestamp 1635444444
transform -1 0 4324 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_42
timestamp 1635444444
transform 1 0 4968 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _222_
timestamp 1635444444
transform 1 0 4692 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_54
timestamp 1635444444
transform 1 0 6072 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1635444444
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1635444444
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1635444444
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1635444444
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_93
timestamp 1635444444
transform 1 0 9660 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_99
timestamp 1635444444
transform 1 0 10212 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1635444444
transform 1 0 9936 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1635444444
transform -1 0 10856 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_90_10
timestamp 1635444444
transform 1 0 2024 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1635444444
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _233_
timestamp 1635444444
transform 1 0 1380 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_90_21
timestamp 1635444444
transform 1 0 3036 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _235_
timestamp 1635444444
transform 1 0 2392 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1635444444
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_90_29
timestamp 1635444444
transform 1 0 3772 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_36
timestamp 1635444444
transform 1 0 4416 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1635444444
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _169_
timestamp 1635444444
transform -1 0 4416 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_48
timestamp 1635444444
transform 1 0 5520 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_60
timestamp 1635444444
transform 1 0 6624 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_72
timestamp 1635444444
transform 1 0 7728 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_85
timestamp 1635444444
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1635444444
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_97
timestamp 1635444444
transform 1 0 10028 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1635444444
transform -1 0 10856 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_10
timestamp 1635444444
transform 1 0 2024 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1635444444
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _232_
timestamp 1635444444
transform 1 0 1380 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_91_18
timestamp 1635444444
transform 1 0 2760 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_25
timestamp 1635444444
transform 1 0 3404 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _221_
timestamp 1635444444
transform 1 0 3128 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1635444444
transform 1 0 2392 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_37
timestamp 1635444444
transform 1 0 4508 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_49
timestamp 1635444444
transform 1 0 5612 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1635444444
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1635444444
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1635444444
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1635444444
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1635444444
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_93
timestamp 1635444444
transform 1 0 9660 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_99
timestamp 1635444444
transform 1 0 10212 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1635444444
transform 1 0 9936 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1635444444
transform -1 0 10856 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_92_7
timestamp 1635444444
transform 1 0 1748 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_7
timestamp 1635444444
transform 1 0 1748 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1635444444
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1635444444
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1635444444
transform -1 0 1748 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1635444444
transform -1 0 1748 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1635444444
transform 1 0 2116 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_13
timestamp 1635444444
transform 1 0 2300 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_17
timestamp 1635444444
transform 1 0 2668 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_24
timestamp 1635444444
transform 1 0 3312 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_15
timestamp 1635444444
transform 1 0 2484 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_22
timestamp 1635444444
transform 1 0 3128 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _223_
timestamp 1635444444
transform 1 0 2392 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _224_
timestamp 1635444444
transform 1 0 3036 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _225_
timestamp 1635444444
transform 1 0 2852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1635444444
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_34
timestamp 1635444444
transform 1 0 4232 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1635444444
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1635444444
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_46
timestamp 1635444444
transform 1 0 5336 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1635444444
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1635444444
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_57
timestamp 1635444444
transform 1 0 6348 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_63
timestamp 1635444444
transform 1 0 6900 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1635444444
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1635444444
transform -1 0 7268 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1635444444
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1635444444
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_67
timestamp 1635444444
transform 1 0 7268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1635444444
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_88
timestamp 1635444444
transform 1 0 9200 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_79
timestamp 1635444444
transform 1 0 8372 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1635444444
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1635444444
transform -1 0 9200 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_99
timestamp 1635444444
transform 1 0 10212 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_91
timestamp 1635444444
transform 1 0 9476 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1635444444
transform 1 0 9936 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1635444444
transform -1 0 10856 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1635444444
transform -1 0 10856 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1635444444
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1635444444
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1635444444
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _231_
timestamp 1635444444
transform 1 0 2024 0 1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_94_20
timestamp 1635444444
transform 1 0 2944 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1635444444
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1635444444
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1635444444
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_53
timestamp 1635444444
transform 1 0 5980 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_57
timestamp 1635444444
transform 1 0 6348 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_62
timestamp 1635444444
transform 1 0 6808 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _175_
timestamp 1635444444
transform -1 0 6808 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_74
timestamp 1635444444
transform 1 0 7912 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_82
timestamp 1635444444
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_85
timestamp 1635444444
transform 1 0 8924 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1635444444
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_94_93
timestamp 1635444444
transform 1 0 9660 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_99
timestamp 1635444444
transform 1 0 10212 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1635444444
transform 1 0 9936 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1635444444
transform -1 0 10856 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_7
timestamp 1635444444
transform 1 0 1748 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1635444444
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1635444444
transform -1 0 1748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_25
timestamp 1635444444
transform 1 0 3404 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _228_
timestamp 1635444444
transform 1 0 2484 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_95_33
timestamp 1635444444
transform 1 0 4140 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _226_
timestamp 1635444444
transform -1 0 4140 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_45
timestamp 1635444444
transform 1 0 5244 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_53
timestamp 1635444444
transform 1 0 5980 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1635444444
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1635444444
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1635444444
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1635444444
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_93
timestamp 1635444444
transform 1 0 9660 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_99
timestamp 1635444444
transform 1 0 10212 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1635444444
transform 1 0 9936 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1635444444
transform -1 0 10856 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_7
timestamp 1635444444
transform 1 0 1748 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1635444444
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1635444444
transform -1 0 1748 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_19
timestamp 1635444444
transform 1 0 2852 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1635444444
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1635444444
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1635444444
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1635444444
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1635444444
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1635444444
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1635444444
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1635444444
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_85
timestamp 1635444444
transform 1 0 8924 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1635444444
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_96_93
timestamp 1635444444
transform 1 0 9660 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_99
timestamp 1635444444
transform 1 0 10212 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1635444444
transform 1 0 9936 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1635444444
transform -1 0 10856 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_10
timestamp 1635444444
transform 1 0 2024 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1635444444
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _243_
timestamp 1635444444
transform 1 0 1380 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_97_18
timestamp 1635444444
transform 1 0 2760 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1635444444
transform 1 0 2392 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_30
timestamp 1635444444
transform 1 0 3864 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_42
timestamp 1635444444
transform 1 0 4968 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_54
timestamp 1635444444
transform 1 0 6072 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1635444444
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1635444444
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1635444444
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1635444444
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_101
timestamp 1635444444
transform 1 0 10396 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_97_93
timestamp 1635444444
transform 1 0 9660 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1635444444
transform -1 0 10856 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_98_3
timestamp 1635444444
transform 1 0 1380 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1635444444
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _238_
timestamp 1635444444
transform 1 0 1932 0 1 55488
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_98_19
timestamp 1635444444
transform 1 0 2852 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1635444444
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_33
timestamp 1635444444
transform 1 0 4140 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1635444444
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1635444444
transform 1 0 3772 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_45
timestamp 1635444444
transform 1 0 5244 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_57
timestamp 1635444444
transform 1 0 6348 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_69
timestamp 1635444444
transform 1 0 7452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_81
timestamp 1635444444
transform 1 0 8556 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_98_85
timestamp 1635444444
transform 1 0 8924 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1635444444
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_93
timestamp 1635444444
transform 1 0 9660 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_99
timestamp 1635444444
transform 1 0 10212 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1635444444
transform 1 0 9844 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1635444444
transform -1 0 10856 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_100_10
timestamp 1635444444
transform 1 0 2024 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_10
timestamp 1635444444
transform 1 0 2024 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1635444444
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1635444444
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _240_
timestamp 1635444444
transform 1 0 1380 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _242_
timestamp 1635444444
transform 1 0 1380 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_100_18
timestamp 1635444444
transform 1 0 2760 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_23
timestamp 1635444444
transform 1 0 3220 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_14
timestamp 1635444444
transform 1 0 2392 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_25
timestamp 1635444444
transform 1 0 3404 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _227_
timestamp 1635444444
transform 1 0 2852 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _237_
timestamp 1635444444
transform 1 0 2484 0 -1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1635444444
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_33
timestamp 1635444444
transform 1 0 4140 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_33
timestamp 1635444444
transform 1 0 4140 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1635444444
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _230_
timestamp 1635444444
transform 1 0 3772 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1635444444
transform 1 0 3772 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_45
timestamp 1635444444
transform 1 0 5244 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_45
timestamp 1635444444
transform 1 0 5244 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_57
timestamp 1635444444
transform 1 0 6348 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_53
timestamp 1635444444
transform 1 0 5980 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1635444444
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1635444444
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_69
timestamp 1635444444
transform 1 0 7452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1635444444
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_81
timestamp 1635444444
transform 1 0 8556 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_85
timestamp 1635444444
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1635444444
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1635444444
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_97
timestamp 1635444444
transform 1 0 10028 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_99_93
timestamp 1635444444
transform 1 0 9660 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_99
timestamp 1635444444
transform 1 0 10212 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1635444444
transform 1 0 9844 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1635444444
transform -1 0 10856 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1635444444
transform -1 0 10856 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_10
timestamp 1635444444
transform 1 0 2024 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1635444444
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _239_
timestamp 1635444444
transform 1 0 1380 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_101_18
timestamp 1635444444
transform 1 0 2760 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1635444444
transform -1 0 2760 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_30
timestamp 1635444444
transform 1 0 3864 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_42
timestamp 1635444444
transform 1 0 4968 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_54
timestamp 1635444444
transform 1 0 6072 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1635444444
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1635444444
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1635444444
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_81
timestamp 1635444444
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_93
timestamp 1635444444
transform 1 0 9660 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_99
timestamp 1635444444
transform 1 0 10212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1635444444
transform 1 0 9844 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1635444444
transform -1 0 10856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_102_10
timestamp 1635444444
transform 1 0 2024 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1635444444
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _241_
timestamp 1635444444
transform 1 0 1380 0 1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_102_18
timestamp 1635444444
transform 1 0 2760 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1635444444
transform 1 0 2392 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_102_26
timestamp 1635444444
transform 1 0 3496 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_102_29
timestamp 1635444444
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1635444444
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_41
timestamp 1635444444
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_53
timestamp 1635444444
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1635444444
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1635444444
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1635444444
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_85
timestamp 1635444444
transform 1 0 8924 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1635444444
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_102_93
timestamp 1635444444
transform 1 0 9660 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_102_99
timestamp 1635444444
transform 1 0 10212 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1635444444
transform 1 0 9844 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1635444444
transform -1 0 10856 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_7
timestamp 1635444444
transform 1 0 1748 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1635444444
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1635444444
transform -1 0 1748 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_19
timestamp 1635444444
transform 1 0 2852 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_31
timestamp 1635444444
transform 1 0 3956 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_43
timestamp 1635444444
transform 1 0 5060 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1635444444
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1635444444
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1635444444
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1635444444
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_81
timestamp 1635444444
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_93
timestamp 1635444444
transform 1 0 9660 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_99
timestamp 1635444444
transform 1 0 10212 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1635444444
transform 1 0 9844 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1635444444
transform -1 0 10856 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_104_7
timestamp 1635444444
transform 1 0 1748 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1635444444
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1635444444
transform -1 0 1748 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_104_19
timestamp 1635444444
transform 1 0 2852 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1635444444
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1635444444
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1635444444
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_41
timestamp 1635444444
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_53
timestamp 1635444444
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_65
timestamp 1635444444
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1635444444
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1635444444
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_85
timestamp 1635444444
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1635444444
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_104_97
timestamp 1635444444
transform 1 0 10028 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1635444444
transform -1 0 10856 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_7
timestamp 1635444444
transform 1 0 1748 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_7
timestamp 1635444444
transform 1 0 1748 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1635444444
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1635444444
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1635444444
transform -1 0 1748 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1635444444
transform -1 0 1748 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_19
timestamp 1635444444
transform 1 0 2852 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_19
timestamp 1635444444
transform 1 0 2852 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_31
timestamp 1635444444
transform 1 0 3956 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1635444444
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1635444444
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1635444444
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_43
timestamp 1635444444
transform 1 0 5060 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1635444444
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1635444444
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1635444444
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1635444444
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1635444444
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1635444444
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_65
timestamp 1635444444
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1635444444
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_105_81
timestamp 1635444444
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1635444444
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_85
timestamp 1635444444
transform 1 0 8924 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1635444444
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_93
timestamp 1635444444
transform 1 0 9660 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_105_99
timestamp 1635444444
transform 1 0 10212 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_93
timestamp 1635444444
transform 1 0 9660 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_99
timestamp 1635444444
transform 1 0 10212 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1635444444
transform 1 0 9844 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1635444444
transform 1 0 9844 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1635444444
transform -1 0 10856 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1635444444
transform -1 0 10856 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_7
timestamp 1635444444
transform 1 0 1748 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1635444444
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1635444444
transform -1 0 1748 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_19
timestamp 1635444444
transform 1 0 2852 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_31
timestamp 1635444444
transform 1 0 3956 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_43
timestamp 1635444444
transform 1 0 5060 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1635444444
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1635444444
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1635444444
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1635444444
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_81
timestamp 1635444444
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_93
timestamp 1635444444
transform 1 0 9660 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_107_99
timestamp 1635444444
transform 1 0 10212 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1635444444
transform 1 0 9844 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1635444444
transform -1 0 10856 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_7
timestamp 1635444444
transform 1 0 1748 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1635444444
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1635444444
transform -1 0 1748 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_19
timestamp 1635444444
transform 1 0 2852 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1635444444
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_29
timestamp 1635444444
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1635444444
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_41
timestamp 1635444444
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_53
timestamp 1635444444
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_65
timestamp 1635444444
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1635444444
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1635444444
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_85
timestamp 1635444444
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1635444444
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_97
timestamp 1635444444
transform 1 0 10028 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1635444444
transform -1 0 10856 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_109_7
timestamp 1635444444
transform 1 0 1748 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1635444444
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1635444444
transform 1 0 2116 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1635444444
transform -1 0 1748 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_109_14
timestamp 1635444444
transform 1 0 2392 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_26
timestamp 1635444444
transform 1 0 3496 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_38
timestamp 1635444444
transform 1 0 4600 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_50
timestamp 1635444444
transform 1 0 5704 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1635444444
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1635444444
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1635444444
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_81
timestamp 1635444444
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_93
timestamp 1635444444
transform 1 0 9660 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_109_99
timestamp 1635444444
transform 1 0 10212 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1635444444
transform 1 0 9844 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1635444444
transform -1 0 10856 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_110_7
timestamp 1635444444
transform 1 0 1748 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1635444444
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1635444444
transform -1 0 1748 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_13
timestamp 1635444444
transform 1 0 2300 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_110_24
timestamp 1635444444
transform 1 0 3312 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _245_
timestamp 1635444444
transform -1 0 3312 0 1 62016
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1635444444
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1635444444
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1635444444
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1635444444
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_65
timestamp 1635444444
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1635444444
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1635444444
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_85
timestamp 1635444444
transform 1 0 8924 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1635444444
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_110_93
timestamp 1635444444
transform 1 0 9660 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_110_99
timestamp 1635444444
transform 1 0 10212 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1635444444
transform 1 0 9844 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1635444444
transform -1 0 10856 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_111_3
timestamp 1635444444
transform 1 0 1380 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1635444444
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _246_
timestamp 1635444444
transform 1 0 1656 0 -1 63104
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_111_13
timestamp 1635444444
transform 1 0 2300 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_17
timestamp 1635444444
transform 1 0 2668 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _244_
timestamp 1635444444
transform 1 0 2760 0 -1 63104
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_111_28
timestamp 1635444444
transform 1 0 3680 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_40
timestamp 1635444444
transform 1 0 4784 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_52
timestamp 1635444444
transform 1 0 5888 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_57
timestamp 1635444444
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1635444444
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_69
timestamp 1635444444
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_81
timestamp 1635444444
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_101
timestamp 1635444444
transform 1 0 10396 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_111_93
timestamp 1635444444
transform 1 0 9660 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1635444444
transform -1 0 10856 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_112_12
timestamp 1635444444
transform 1 0 2208 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_112_3
timestamp 1635444444
transform 1 0 1380 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_113_11
timestamp 1635444444
transform 1 0 2116 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_3
timestamp 1635444444
transform 1 0 1380 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1635444444
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1635444444
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _247_
timestamp 1635444444
transform 1 0 1564 0 1 63104
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _248_
timestamp 1635444444
transform 1 0 1472 0 -1 64192
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_112_19
timestamp 1635444444
transform 1 0 2852 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_22
timestamp 1635444444
transform 1 0 3128 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _250_
timestamp 1635444444
transform 1 0 2484 0 -1 64192
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1635444444
transform 1 0 2576 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1635444444
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_32
timestamp 1635444444
transform 1 0 4048 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_34
timestamp 1635444444
transform 1 0 4232 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1635444444
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1635444444
transform 1 0 3772 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_44
timestamp 1635444444
transform 1 0 5152 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_46
timestamp 1635444444
transform 1 0 5336 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_56
timestamp 1635444444
transform 1 0 6256 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_54
timestamp 1635444444
transform 1 0 6072 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1635444444
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1635444444
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_68
timestamp 1635444444
transform 1 0 7360 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1635444444
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_112_80
timestamp 1635444444
transform 1 0 8464 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_112_85
timestamp 1635444444
transform 1 0 8924 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_81
timestamp 1635444444
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1635444444
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_112_93
timestamp 1635444444
transform 1 0 9660 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_112_99
timestamp 1635444444
transform 1 0 10212 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_113_93
timestamp 1635444444
transform 1 0 9660 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_113_99
timestamp 1635444444
transform 1 0 10212 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1635444444
transform 1 0 9844 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1635444444
transform 1 0 9844 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1635444444
transform -1 0 10856 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1635444444
transform -1 0 10856 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_114_11
timestamp 1635444444
transform 1 0 2116 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_114_3
timestamp 1635444444
transform 1 0 1380 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1635444444
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _249_
timestamp 1635444444
transform 1 0 1472 0 1 64192
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_114_18
timestamp 1635444444
transform 1 0 2760 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1635444444
transform 1 0 2484 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_114_26
timestamp 1635444444
transform 1 0 3496 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_114_29
timestamp 1635444444
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1635444444
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_41
timestamp 1635444444
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_53
timestamp 1635444444
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_65
timestamp 1635444444
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1635444444
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1635444444
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_85
timestamp 1635444444
transform 1 0 8924 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1635444444
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_114_93
timestamp 1635444444
transform 1 0 9660 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_114_99
timestamp 1635444444
transform 1 0 10212 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1635444444
transform 1 0 9844 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1635444444
transform -1 0 10856 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_115_6
timestamp 1635444444
transform 1 0 1656 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1635444444
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1635444444
transform -1 0 1656 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_21
timestamp 1635444444
transform 1 0 3036 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _253_
timestamp 1635444444
transform 1 0 2392 0 -1 65280
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_115_33
timestamp 1635444444
transform 1 0 4140 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_45
timestamp 1635444444
transform 1 0 5244 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_115_53
timestamp 1635444444
transform 1 0 5980 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_57
timestamp 1635444444
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1635444444
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_69
timestamp 1635444444
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_81
timestamp 1635444444
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_115_101
timestamp 1635444444
transform 1 0 10396 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_115_93
timestamp 1635444444
transform 1 0 9660 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1635444444
transform -1 0 10856 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_116_6
timestamp 1635444444
transform 1 0 1656 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1635444444
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1635444444
transform -1 0 1656 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_116_24
timestamp 1635444444
transform 1 0 3312 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _252_
timestamp 1635444444
transform -1 0 3312 0 1 65280
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1635444444
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _251_
timestamp 1635444444
transform 1 0 3772 0 1 65280
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_116_39
timestamp 1635444444
transform 1 0 4692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_51
timestamp 1635444444
transform 1 0 5796 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_63
timestamp 1635444444
transform 1 0 6900 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_75
timestamp 1635444444
transform 1 0 8004 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1635444444
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_85
timestamp 1635444444
transform 1 0 8924 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1635444444
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_116_93
timestamp 1635444444
transform 1 0 9660 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_116_99
timestamp 1635444444
transform 1 0 10212 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1635444444
transform 1 0 9844 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1635444444
transform -1 0 10856 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_10
timestamp 1635444444
transform 1 0 2024 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1635444444
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _257_
timestamp 1635444444
transform 1 0 1380 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_117_21
timestamp 1635444444
transform 1 0 3036 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _254_
timestamp 1635444444
transform 1 0 2392 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _256_
timestamp 1635444444
transform 1 0 3404 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_117_32
timestamp 1635444444
transform 1 0 4048 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_44
timestamp 1635444444
transform 1 0 5152 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1635444444
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1635444444
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1635444444
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_81
timestamp 1635444444
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_117_93
timestamp 1635444444
transform 1 0 9660 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_117_99
timestamp 1635444444
transform 1 0 10212 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1635444444
transform 1 0 9844 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1635444444
transform -1 0 10856 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_118_6
timestamp 1635444444
transform 1 0 1656 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_119_6
timestamp 1635444444
transform 1 0 1656 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1635444444
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1635444444
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1635444444
transform -1 0 1656 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1635444444
transform -1 0 1656 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1635444444
transform 1 0 2024 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_118_21
timestamp 1635444444
transform 1 0 3036 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_119_13
timestamp 1635444444
transform 1 0 2300 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_25
timestamp 1635444444
transform 1 0 3404 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _255_
timestamp 1635444444
transform 1 0 2392 0 1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1635444444
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_29
timestamp 1635444444
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_37
timestamp 1635444444
transform 1 0 4508 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1635444444
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_41
timestamp 1635444444
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_49
timestamp 1635444444
transform 1 0 5612 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_118_53
timestamp 1635444444
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1635444444
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1635444444
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1635444444
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_65
timestamp 1635444444
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1635444444
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_119_69
timestamp 1635444444
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1635444444
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_85
timestamp 1635444444
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_81
timestamp 1635444444
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1635444444
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_118_97
timestamp 1635444444
transform 1 0 10028 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_119_93
timestamp 1635444444
transform 1 0 9660 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_119_99
timestamp 1635444444
transform 1 0 10212 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1635444444
transform 1 0 9844 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1635444444
transform -1 0 10856 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1635444444
transform -1 0 10856 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_6
timestamp 1635444444
transform 1 0 1656 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1635444444
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1635444444
transform -1 0 1656 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1635444444
transform 1 0 2024 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_120_13
timestamp 1635444444
transform 1 0 2300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_25
timestamp 1635444444
transform 1 0 3404 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_120_29
timestamp 1635444444
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1635444444
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_41
timestamp 1635444444
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_53
timestamp 1635444444
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_65
timestamp 1635444444
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1635444444
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1635444444
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_85
timestamp 1635444444
transform 1 0 8924 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1635444444
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_120_93
timestamp 1635444444
transform 1 0 9660 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_120_99
timestamp 1635444444
transform 1 0 10212 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1635444444
transform 1 0 9844 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1635444444
transform -1 0 10856 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_121_6
timestamp 1635444444
transform 1 0 1656 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1635444444
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1635444444
transform -1 0 1656 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_121_18
timestamp 1635444444
transform 1 0 2760 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_30
timestamp 1635444444
transform 1 0 3864 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_42
timestamp 1635444444
transform 1 0 4968 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_54
timestamp 1635444444
transform 1 0 6072 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1635444444
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1635444444
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1635444444
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_81
timestamp 1635444444
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_93
timestamp 1635444444
transform 1 0 9660 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_121_99
timestamp 1635444444
transform 1 0 10212 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1635444444
transform 1 0 9844 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1635444444
transform -1 0 10856 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_122_6
timestamp 1635444444
transform 1 0 1656 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1635444444
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1635444444
transform -1 0 1656 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_122_18
timestamp 1635444444
transform 1 0 2760 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_122_26
timestamp 1635444444
transform 1 0 3496 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_122_29
timestamp 1635444444
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1635444444
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_41
timestamp 1635444444
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_53
timestamp 1635444444
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_65
timestamp 1635444444
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1635444444
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1635444444
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_85
timestamp 1635444444
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1635444444
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_122_97
timestamp 1635444444
transform 1 0 10028 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1635444444
transform -1 0 10856 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_6
timestamp 1635444444
transform 1 0 1656 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1635444444
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1635444444
transform -1 0 1656 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_18
timestamp 1635444444
transform 1 0 2760 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_30
timestamp 1635444444
transform 1 0 3864 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_42
timestamp 1635444444
transform 1 0 4968 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_54
timestamp 1635444444
transform 1 0 6072 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_57
timestamp 1635444444
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1635444444
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_69
timestamp 1635444444
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_81
timestamp 1635444444
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_93
timestamp 1635444444
transform 1 0 9660 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_123_99
timestamp 1635444444
transform 1 0 10212 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1635444444
transform 1 0 9844 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1635444444
transform -1 0 10856 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_124_6
timestamp 1635444444
transform 1 0 1656 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1635444444
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1635444444
transform -1 0 1656 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_124_18
timestamp 1635444444
transform 1 0 2760 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_124_26
timestamp 1635444444
transform 1 0 3496 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_124_29
timestamp 1635444444
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1635444444
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_41
timestamp 1635444444
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_53
timestamp 1635444444
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_65
timestamp 1635444444
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1635444444
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1635444444
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_85
timestamp 1635444444
transform 1 0 8924 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1635444444
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_124_93
timestamp 1635444444
transform 1 0 9660 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_124_99
timestamp 1635444444
transform 1 0 10212 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1635444444
transform 1 0 9844 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1635444444
transform -1 0 10856 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_6
timestamp 1635444444
transform 1 0 1656 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_6
timestamp 1635444444
transform 1 0 1656 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1635444444
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1635444444
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1635444444
transform -1 0 1656 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1635444444
transform -1 0 1656 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_18
timestamp 1635444444
transform 1 0 2760 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_18
timestamp 1635444444
transform 1 0 2760 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_125_30
timestamp 1635444444
transform 1 0 3864 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_126_26
timestamp 1635444444
transform 1 0 3496 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1635444444
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _259_
timestamp 1635444444
transform 1 0 3772 0 1 70720
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_125_42
timestamp 1635444444
transform 1 0 4968 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_39
timestamp 1635444444
transform 1 0 4692 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_51
timestamp 1635444444
transform 1 0 5796 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_125_54
timestamp 1635444444
transform 1 0 6072 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_125_57
timestamp 1635444444
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_63
timestamp 1635444444
transform 1 0 6900 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1635444444
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_69
timestamp 1635444444
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_75
timestamp 1635444444
transform 1 0 8004 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_125_81
timestamp 1635444444
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1635444444
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_85
timestamp 1635444444
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1635444444
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_125_93
timestamp 1635444444
transform 1 0 9660 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_125_99
timestamp 1635444444
transform 1 0 10212 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_126_97
timestamp 1635444444
transform 1 0 10028 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1635444444
transform 1 0 9844 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1635444444
transform -1 0 10856 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1635444444
transform -1 0 10856 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_6
timestamp 1635444444
transform 1 0 1656 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1635444444
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _260_
timestamp 1635444444
transform 1 0 2024 0 -1 71808
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1635444444
transform -1 0 1656 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_17
timestamp 1635444444
transform 1 0 2668 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _258_
timestamp 1635444444
transform -1 0 3956 0 -1 71808
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_127_31
timestamp 1635444444
transform 1 0 3956 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_43
timestamp 1635444444
transform 1 0 5060 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1635444444
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_57
timestamp 1635444444
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1635444444
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_69
timestamp 1635444444
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_81
timestamp 1635444444
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_93
timestamp 1635444444
transform 1 0 9660 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_127_99
timestamp 1635444444
transform 1 0 10212 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1635444444
transform 1 0 9844 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1635444444
transform -1 0 10856 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_128_6
timestamp 1635444444
transform 1 0 1656 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1635444444
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1635444444
transform -1 0 1656 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_128_14
timestamp 1635444444
transform 1 0 2392 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_128_22
timestamp 1635444444
transform 1 0 3128 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _261_
timestamp 1635444444
transform 1 0 2484 0 1 71808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_128_36
timestamp 1635444444
transform 1 0 4416 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1635444444
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _262_
timestamp 1635444444
transform 1 0 3772 0 1 71808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_128_48
timestamp 1635444444
transform 1 0 5520 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_60
timestamp 1635444444
transform 1 0 6624 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_72
timestamp 1635444444
transform 1 0 7728 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_85
timestamp 1635444444
transform 1 0 8924 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1635444444
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_128_93
timestamp 1635444444
transform 1 0 9660 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_128_99
timestamp 1635444444
transform 1 0 10212 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1635444444
transform 1 0 9844 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1635444444
transform -1 0 10856 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_129_6
timestamp 1635444444
transform 1 0 1656 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1635444444
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1635444444
transform -1 0 1656 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1635444444
transform -1 0 2300 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_129_13
timestamp 1635444444
transform 1 0 2300 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _265_
timestamp 1635444444
transform 1 0 2668 0 -1 72896
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_129_27
timestamp 1635444444
transform 1 0 3588 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _266_
timestamp 1635444444
transform 1 0 3956 0 -1 72896
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_129_41
timestamp 1635444444
transform 1 0 4876 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_129_53
timestamp 1635444444
transform 1 0 5980 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_129_57
timestamp 1635444444
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1635444444
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_69
timestamp 1635444444
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_81
timestamp 1635444444
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_101
timestamp 1635444444
transform 1 0 10396 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_129_93
timestamp 1635444444
transform 1 0 9660 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1635444444
transform -1 0 10856 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_130_10
timestamp 1635444444
transform 1 0 2024 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1635444444
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _271_
timestamp 1635444444
transform 1 0 1380 0 1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_130_14
timestamp 1635444444
transform 1 0 2392 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_130_22
timestamp 1635444444
transform 1 0 3128 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _263_
timestamp 1635444444
transform 1 0 2484 0 1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_130_29
timestamp 1635444444
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1635444444
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_41
timestamp 1635444444
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_53
timestamp 1635444444
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_65
timestamp 1635444444
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1635444444
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1635444444
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_85
timestamp 1635444444
transform 1 0 8924 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1635444444
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_130_93
timestamp 1635444444
transform 1 0 9660 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_130_99
timestamp 1635444444
transform 1 0 10212 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1635444444
transform 1 0 9844 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1635444444
transform -1 0 10856 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_131_10
timestamp 1635444444
transform 1 0 2024 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1635444444
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _267_
timestamp 1635444444
transform 1 0 1380 0 -1 73984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_131_14
timestamp 1635444444
transform 1 0 2392 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_131_22
timestamp 1635444444
transform 1 0 3128 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _264_
timestamp 1635444444
transform 1 0 2484 0 -1 73984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_131_33
timestamp 1635444444
transform 1 0 4140 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _273_
timestamp 1635444444
transform 1 0 3496 0 -1 73984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _274_
timestamp 1635444444
transform 1 0 4508 0 -1 73984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_131_44
timestamp 1635444444
transform 1 0 5152 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_57
timestamp 1635444444
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1635444444
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_69
timestamp 1635444444
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_81
timestamp 1635444444
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_93
timestamp 1635444444
transform 1 0 9660 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_131_99
timestamp 1635444444
transform 1 0 10212 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1635444444
transform 1 0 9844 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1635444444
transform -1 0 10856 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_10
timestamp 1635444444
transform 1 0 2024 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_133_10
timestamp 1635444444
transform 1 0 2024 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1635444444
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1635444444
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _268_
timestamp 1635444444
transform 1 0 1380 0 1 73984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _269_
timestamp 1635444444
transform 1 0 1380 0 -1 75072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_132_21
timestamp 1635444444
transform 1 0 3036 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_133_21
timestamp 1635444444
transform 1 0 3036 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _270_
timestamp 1635444444
transform 1 0 2392 0 1 73984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _272_
timestamp 1635444444
transform 1 0 2392 0 -1 75072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1635444444
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_32
timestamp 1635444444
transform 1 0 4048 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_33
timestamp 1635444444
transform 1 0 4140 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1635444444
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1635444444
transform -1 0 4048 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_44
timestamp 1635444444
transform 1 0 5152 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_45
timestamp 1635444444
transform 1 0 5244 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_132_56
timestamp 1635444444
transform 1 0 6256 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_133_53
timestamp 1635444444
transform 1 0 5980 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_133_57
timestamp 1635444444
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1635444444
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_68
timestamp 1635444444
transform 1 0 7360 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_69
timestamp 1635444444
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_132_80
timestamp 1635444444
transform 1 0 8464 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_132_85
timestamp 1635444444
transform 1 0 8924 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_81
timestamp 1635444444
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1635444444
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_132_93
timestamp 1635444444
transform 1 0 9660 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_132_99
timestamp 1635444444
transform 1 0 10212 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_133_101
timestamp 1635444444
transform 1 0 10396 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_133_93
timestamp 1635444444
transform 1 0 9660 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1635444444
transform 1 0 9844 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1635444444
transform -1 0 10856 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1635444444
transform -1 0 10856 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_6
timestamp 1635444444
transform 1 0 1656 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1635444444
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1635444444
transform -1 0 1656 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1635444444
transform -1 0 2300 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_134_13
timestamp 1635444444
transform 1 0 2300 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_134_25
timestamp 1635444444
transform 1 0 3404 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_134_29
timestamp 1635444444
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1635444444
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_41
timestamp 1635444444
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_53
timestamp 1635444444
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_65
timestamp 1635444444
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1635444444
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1635444444
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_85
timestamp 1635444444
transform 1 0 8924 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1635444444
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_134_93
timestamp 1635444444
transform 1 0 9660 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_134_99
timestamp 1635444444
transform 1 0 10212 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1635444444
transform 1 0 9844 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1635444444
transform -1 0 10856 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_6
timestamp 1635444444
transform 1 0 1656 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1635444444
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1635444444
transform -1 0 1656 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_18
timestamp 1635444444
transform 1 0 2760 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_30
timestamp 1635444444
transform 1 0 3864 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_42
timestamp 1635444444
transform 1 0 4968 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_135_54
timestamp 1635444444
transform 1 0 6072 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_135_57
timestamp 1635444444
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1635444444
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_69
timestamp 1635444444
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_81
timestamp 1635444444
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_135_93
timestamp 1635444444
transform 1 0 9660 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_135_99
timestamp 1635444444
transform 1 0 10212 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1635444444
transform 1 0 9844 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1635444444
transform -1 0 10856 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_136_6
timestamp 1635444444
transform 1 0 1656 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1635444444
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1635444444
transform -1 0 1656 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_136_18
timestamp 1635444444
transform 1 0 2760 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_136_26
timestamp 1635444444
transform 1 0 3496 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_136_29
timestamp 1635444444
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1635444444
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_41
timestamp 1635444444
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_53
timestamp 1635444444
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_65
timestamp 1635444444
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1635444444
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1635444444
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_85
timestamp 1635444444
transform 1 0 8924 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1635444444
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_136_93
timestamp 1635444444
transform 1 0 9660 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_136_99
timestamp 1635444444
transform 1 0 10212 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1635444444
transform 1 0 9844 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1635444444
transform -1 0 10856 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_6
timestamp 1635444444
transform 1 0 1656 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1635444444
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1635444444
transform -1 0 1656 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1635444444
transform -1 0 2300 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_13
timestamp 1635444444
transform 1 0 2300 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_137_20
timestamp 1635444444
transform 1 0 2944 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1635444444
transform -1 0 2944 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_137_32
timestamp 1635444444
transform 1 0 4048 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_44
timestamp 1635444444
transform 1 0 5152 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_57
timestamp 1635444444
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1635444444
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_69
timestamp 1635444444
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_81
timestamp 1635444444
transform 1 0 8556 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1635444444
transform 1 0 9108 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_91
timestamp 1635444444
transform 1 0 9476 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_99
timestamp 1635444444
transform 1 0 10212 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1635444444
transform 1 0 9844 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1635444444
transform -1 0 10856 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_6
timestamp 1635444444
transform 1 0 1656 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1635444444
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1635444444
transform -1 0 1656 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1635444444
transform -1 0 2300 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_13
timestamp 1635444444
transform 1 0 2300 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_138_20
timestamp 1635444444
transform 1 0 2944 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1635444444
transform 1 0 2668 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_32
timestamp 1635444444
transform 1 0 4048 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1635444444
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1635444444
transform -1 0 4048 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_44
timestamp 1635444444
transform 1 0 5152 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_57
timestamp 1635444444
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1635444444
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_69
timestamp 1635444444
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1635444444
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_138_85
timestamp 1635444444
transform 1 0 8924 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1635444444
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1635444444
transform 1 0 9108 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_91
timestamp 1635444444
transform 1 0 9476 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_99
timestamp 1635444444
transform 1 0 10212 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1635444444
transform 1 0 9844 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1635444444
transform -1 0 10856 0 1 77248
box -38 -48 314 592
<< labels >>
rlabel metal4 s 2575 2128 2895 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 5839 2128 6159 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 9103 2128 9423 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 4207 2128 4527 77840 6 vssd1
port 1 nsew ground input
rlabel metal4 s 7471 2128 7791 77840 6 vssd1
port 1 nsew ground input
rlabel metal3 s 11200 280 12000 400 6 wb_clk_i
port 2 nsew signal input
rlabel metal3 s 11200 960 12000 1080 6 wb_rst_i
port 3 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wbs_hr_ack_i
port 4 nsew signal input
rlabel metal3 s 0 824 800 944 6 wbs_hr_cyc_o
port 5 nsew signal tristate
rlabel metal3 s 0 22448 800 22568 6 wbs_hr_dat_i[0]
port 6 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 wbs_hr_dat_i[10]
port 7 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 wbs_hr_dat_i[11]
port 8 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 wbs_hr_dat_i[12]
port 9 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 wbs_hr_dat_i[13]
port 10 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 wbs_hr_dat_i[14]
port 11 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 wbs_hr_dat_i[15]
port 12 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 wbs_hr_dat_i[16]
port 13 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 wbs_hr_dat_i[17]
port 14 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 wbs_hr_dat_i[18]
port 15 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wbs_hr_dat_i[19]
port 16 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 wbs_hr_dat_i[1]
port 17 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 wbs_hr_dat_i[20]
port 18 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wbs_hr_dat_i[21]
port 19 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 wbs_hr_dat_i[22]
port 20 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 wbs_hr_dat_i[23]
port 21 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 wbs_hr_dat_i[24]
port 22 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 wbs_hr_dat_i[25]
port 23 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 wbs_hr_dat_i[26]
port 24 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 wbs_hr_dat_i[27]
port 25 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 wbs_hr_dat_i[28]
port 26 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 wbs_hr_dat_i[29]
port 27 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 wbs_hr_dat_i[2]
port 28 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 wbs_hr_dat_i[30]
port 29 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 wbs_hr_dat_i[31]
port 30 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 wbs_hr_dat_i[3]
port 31 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 wbs_hr_dat_i[4]
port 32 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wbs_hr_dat_i[5]
port 33 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wbs_hr_dat_i[6]
port 34 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 wbs_hr_dat_i[7]
port 35 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 wbs_hr_dat_i[8]
port 36 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 wbs_hr_dat_i[9]
port 37 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 wbs_hr_dat_o[0]
port 38 nsew signal tristate
rlabel metal3 s 0 9664 800 9784 6 wbs_hr_dat_o[10]
port 39 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 wbs_hr_dat_o[11]
port 40 nsew signal tristate
rlabel metal3 s 0 10752 800 10872 6 wbs_hr_dat_o[12]
port 41 nsew signal tristate
rlabel metal3 s 0 11296 800 11416 6 wbs_hr_dat_o[13]
port 42 nsew signal tristate
rlabel metal3 s 0 11840 800 11960 6 wbs_hr_dat_o[14]
port 43 nsew signal tristate
rlabel metal3 s 0 12384 800 12504 6 wbs_hr_dat_o[15]
port 44 nsew signal tristate
rlabel metal3 s 0 12928 800 13048 6 wbs_hr_dat_o[16]
port 45 nsew signal tristate
rlabel metal3 s 0 13608 800 13728 6 wbs_hr_dat_o[17]
port 46 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 wbs_hr_dat_o[18]
port 47 nsew signal tristate
rlabel metal3 s 0 14696 800 14816 6 wbs_hr_dat_o[19]
port 48 nsew signal tristate
rlabel metal3 s 0 4632 800 4752 6 wbs_hr_dat_o[1]
port 49 nsew signal tristate
rlabel metal3 s 0 15240 800 15360 6 wbs_hr_dat_o[20]
port 50 nsew signal tristate
rlabel metal3 s 0 15784 800 15904 6 wbs_hr_dat_o[21]
port 51 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 wbs_hr_dat_o[22]
port 52 nsew signal tristate
rlabel metal3 s 0 16872 800 16992 6 wbs_hr_dat_o[23]
port 53 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 wbs_hr_dat_o[24]
port 54 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 wbs_hr_dat_o[25]
port 55 nsew signal tristate
rlabel metal3 s 0 18504 800 18624 6 wbs_hr_dat_o[26]
port 56 nsew signal tristate
rlabel metal3 s 0 19048 800 19168 6 wbs_hr_dat_o[27]
port 57 nsew signal tristate
rlabel metal3 s 0 19592 800 19712 6 wbs_hr_dat_o[28]
port 58 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 wbs_hr_dat_o[29]
port 59 nsew signal tristate
rlabel metal3 s 0 5176 800 5296 6 wbs_hr_dat_o[2]
port 60 nsew signal tristate
rlabel metal3 s 0 20816 800 20936 6 wbs_hr_dat_o[30]
port 61 nsew signal tristate
rlabel metal3 s 0 21360 800 21480 6 wbs_hr_dat_o[31]
port 62 nsew signal tristate
rlabel metal3 s 0 5720 800 5840 6 wbs_hr_dat_o[3]
port 63 nsew signal tristate
rlabel metal3 s 0 6264 800 6384 6 wbs_hr_dat_o[4]
port 64 nsew signal tristate
rlabel metal3 s 0 6944 800 7064 6 wbs_hr_dat_o[5]
port 65 nsew signal tristate
rlabel metal3 s 0 7488 800 7608 6 wbs_hr_dat_o[6]
port 66 nsew signal tristate
rlabel metal3 s 0 8032 800 8152 6 wbs_hr_dat_o[7]
port 67 nsew signal tristate
rlabel metal3 s 0 8576 800 8696 6 wbs_hr_dat_o[8]
port 68 nsew signal tristate
rlabel metal3 s 0 9120 800 9240 6 wbs_hr_dat_o[9]
port 69 nsew signal tristate
rlabel metal3 s 0 1912 800 2032 6 wbs_hr_sel_o[0]
port 70 nsew signal tristate
rlabel metal3 s 0 2456 800 2576 6 wbs_hr_sel_o[1]
port 71 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 wbs_hr_sel_o[2]
port 72 nsew signal tristate
rlabel metal3 s 0 3544 800 3664 6 wbs_hr_sel_o[3]
port 73 nsew signal tristate
rlabel metal3 s 0 280 800 400 6 wbs_hr_stb_o
port 74 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 wbs_hr_we_o
port 75 nsew signal tristate
rlabel metal3 s 0 61888 800 62008 6 wbs_or_ack_i
port 76 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 wbs_or_cyc_o
port 77 nsew signal tristate
rlabel metal3 s 0 62432 800 62552 6 wbs_or_dat_i[0]
port 78 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 wbs_or_dat_i[10]
port 79 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 wbs_or_dat_i[11]
port 80 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 wbs_or_dat_i[12]
port 81 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 wbs_or_dat_i[13]
port 82 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 wbs_or_dat_i[14]
port 83 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 wbs_or_dat_i[15]
port 84 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 wbs_or_dat_i[16]
port 85 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 wbs_or_dat_i[17]
port 86 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 wbs_or_dat_i[18]
port 87 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 wbs_or_dat_i[19]
port 88 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 wbs_or_dat_i[1]
port 89 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 wbs_or_dat_i[20]
port 90 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 wbs_or_dat_i[21]
port 91 nsew signal input
rlabel metal3 s 0 74672 800 74792 6 wbs_or_dat_i[22]
port 92 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 wbs_or_dat_i[23]
port 93 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 wbs_or_dat_i[24]
port 94 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 wbs_or_dat_i[25]
port 95 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 wbs_or_dat_i[26]
port 96 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 wbs_or_dat_i[27]
port 97 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 wbs_or_dat_i[28]
port 98 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 wbs_or_dat_i[29]
port 99 nsew signal input
rlabel metal3 s 0 63520 800 63640 6 wbs_or_dat_i[2]
port 100 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 wbs_or_dat_i[30]
port 101 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 wbs_or_dat_i[31]
port 102 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 wbs_or_dat_i[3]
port 103 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 wbs_or_dat_i[4]
port 104 nsew signal input
rlabel metal3 s 0 65152 800 65272 6 wbs_or_dat_i[5]
port 105 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 wbs_or_dat_i[6]
port 106 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 wbs_or_dat_i[7]
port 107 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 wbs_or_dat_i[8]
port 108 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 wbs_or_dat_i[9]
port 109 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 wbs_or_dat_o[0]
port 110 nsew signal tristate
rlabel metal3 s 0 49648 800 49768 6 wbs_or_dat_o[10]
port 111 nsew signal tristate
rlabel metal3 s 0 50192 800 50312 6 wbs_or_dat_o[11]
port 112 nsew signal tristate
rlabel metal3 s 0 50736 800 50856 6 wbs_or_dat_o[12]
port 113 nsew signal tristate
rlabel metal3 s 0 51280 800 51400 6 wbs_or_dat_o[13]
port 114 nsew signal tristate
rlabel metal3 s 0 51824 800 51944 6 wbs_or_dat_o[14]
port 115 nsew signal tristate
rlabel metal3 s 0 52368 800 52488 6 wbs_or_dat_o[15]
port 116 nsew signal tristate
rlabel metal3 s 0 52912 800 53032 6 wbs_or_dat_o[16]
port 117 nsew signal tristate
rlabel metal3 s 0 53592 800 53712 6 wbs_or_dat_o[17]
port 118 nsew signal tristate
rlabel metal3 s 0 54136 800 54256 6 wbs_or_dat_o[18]
port 119 nsew signal tristate
rlabel metal3 s 0 54680 800 54800 6 wbs_or_dat_o[19]
port 120 nsew signal tristate
rlabel metal3 s 0 44616 800 44736 6 wbs_or_dat_o[1]
port 121 nsew signal tristate
rlabel metal3 s 0 55224 800 55344 6 wbs_or_dat_o[20]
port 122 nsew signal tristate
rlabel metal3 s 0 55768 800 55888 6 wbs_or_dat_o[21]
port 123 nsew signal tristate
rlabel metal3 s 0 56312 800 56432 6 wbs_or_dat_o[22]
port 124 nsew signal tristate
rlabel metal3 s 0 56856 800 56976 6 wbs_or_dat_o[23]
port 125 nsew signal tristate
rlabel metal3 s 0 57400 800 57520 6 wbs_or_dat_o[24]
port 126 nsew signal tristate
rlabel metal3 s 0 57944 800 58064 6 wbs_or_dat_o[25]
port 127 nsew signal tristate
rlabel metal3 s 0 58488 800 58608 6 wbs_or_dat_o[26]
port 128 nsew signal tristate
rlabel metal3 s 0 59032 800 59152 6 wbs_or_dat_o[27]
port 129 nsew signal tristate
rlabel metal3 s 0 59576 800 59696 6 wbs_or_dat_o[28]
port 130 nsew signal tristate
rlabel metal3 s 0 60256 800 60376 6 wbs_or_dat_o[29]
port 131 nsew signal tristate
rlabel metal3 s 0 45160 800 45280 6 wbs_or_dat_o[2]
port 132 nsew signal tristate
rlabel metal3 s 0 60800 800 60920 6 wbs_or_dat_o[30]
port 133 nsew signal tristate
rlabel metal3 s 0 61344 800 61464 6 wbs_or_dat_o[31]
port 134 nsew signal tristate
rlabel metal3 s 0 45704 800 45824 6 wbs_or_dat_o[3]
port 135 nsew signal tristate
rlabel metal3 s 0 46248 800 46368 6 wbs_or_dat_o[4]
port 136 nsew signal tristate
rlabel metal3 s 0 46928 800 47048 6 wbs_or_dat_o[5]
port 137 nsew signal tristate
rlabel metal3 s 0 47472 800 47592 6 wbs_or_dat_o[6]
port 138 nsew signal tristate
rlabel metal3 s 0 48016 800 48136 6 wbs_or_dat_o[7]
port 139 nsew signal tristate
rlabel metal3 s 0 48560 800 48680 6 wbs_or_dat_o[8]
port 140 nsew signal tristate
rlabel metal3 s 0 49104 800 49224 6 wbs_or_dat_o[9]
port 141 nsew signal tristate
rlabel metal3 s 0 41896 800 42016 6 wbs_or_sel_o[0]
port 142 nsew signal tristate
rlabel metal3 s 0 42440 800 42560 6 wbs_or_sel_o[1]
port 143 nsew signal tristate
rlabel metal3 s 0 42984 800 43104 6 wbs_or_sel_o[2]
port 144 nsew signal tristate
rlabel metal3 s 0 43528 800 43648 6 wbs_or_sel_o[3]
port 145 nsew signal tristate
rlabel metal3 s 0 40264 800 40384 6 wbs_or_stb_o
port 146 nsew signal tristate
rlabel metal3 s 0 41352 800 41472 6 wbs_or_we_o
port 147 nsew signal tristate
rlabel metal3 s 11200 55224 12000 55344 6 wbs_ufp_ack_o
port 148 nsew signal tristate
rlabel metal3 s 11200 6944 12000 7064 6 wbs_ufp_adr_i[0]
port 149 nsew signal input
rlabel metal3 s 11200 14560 12000 14680 6 wbs_ufp_adr_i[10]
port 150 nsew signal input
rlabel metal3 s 11200 15240 12000 15360 6 wbs_ufp_adr_i[11]
port 151 nsew signal input
rlabel metal3 s 11200 16056 12000 16176 6 wbs_ufp_adr_i[12]
port 152 nsew signal input
rlabel metal3 s 11200 16872 12000 16992 6 wbs_ufp_adr_i[13]
port 153 nsew signal input
rlabel metal3 s 11200 17552 12000 17672 6 wbs_ufp_adr_i[14]
port 154 nsew signal input
rlabel metal3 s 11200 18368 12000 18488 6 wbs_ufp_adr_i[15]
port 155 nsew signal input
rlabel metal3 s 11200 19048 12000 19168 6 wbs_ufp_adr_i[16]
port 156 nsew signal input
rlabel metal3 s 11200 19864 12000 19984 6 wbs_ufp_adr_i[17]
port 157 nsew signal input
rlabel metal3 s 11200 20544 12000 20664 6 wbs_ufp_adr_i[18]
port 158 nsew signal input
rlabel metal3 s 11200 21360 12000 21480 6 wbs_ufp_adr_i[19]
port 159 nsew signal input
rlabel metal3 s 11200 7760 12000 7880 6 wbs_ufp_adr_i[1]
port 160 nsew signal input
rlabel metal3 s 11200 22040 12000 22160 6 wbs_ufp_adr_i[20]
port 161 nsew signal input
rlabel metal3 s 11200 22856 12000 22976 6 wbs_ufp_adr_i[21]
port 162 nsew signal input
rlabel metal3 s 11200 23536 12000 23656 6 wbs_ufp_adr_i[22]
port 163 nsew signal input
rlabel metal3 s 11200 24352 12000 24472 6 wbs_ufp_adr_i[23]
port 164 nsew signal input
rlabel metal3 s 11200 25168 12000 25288 6 wbs_ufp_adr_i[24]
port 165 nsew signal input
rlabel metal3 s 11200 25848 12000 25968 6 wbs_ufp_adr_i[25]
port 166 nsew signal input
rlabel metal3 s 11200 26664 12000 26784 6 wbs_ufp_adr_i[26]
port 167 nsew signal input
rlabel metal3 s 11200 27344 12000 27464 6 wbs_ufp_adr_i[27]
port 168 nsew signal input
rlabel metal3 s 11200 28160 12000 28280 6 wbs_ufp_adr_i[28]
port 169 nsew signal input
rlabel metal3 s 11200 28840 12000 28960 6 wbs_ufp_adr_i[29]
port 170 nsew signal input
rlabel metal3 s 11200 8576 12000 8696 6 wbs_ufp_adr_i[2]
port 171 nsew signal input
rlabel metal3 s 11200 29656 12000 29776 6 wbs_ufp_adr_i[30]
port 172 nsew signal input
rlabel metal3 s 11200 30336 12000 30456 6 wbs_ufp_adr_i[31]
port 173 nsew signal input
rlabel metal3 s 11200 9256 12000 9376 6 wbs_ufp_adr_i[3]
port 174 nsew signal input
rlabel metal3 s 11200 10072 12000 10192 6 wbs_ufp_adr_i[4]
port 175 nsew signal input
rlabel metal3 s 11200 10752 12000 10872 6 wbs_ufp_adr_i[5]
port 176 nsew signal input
rlabel metal3 s 11200 11568 12000 11688 6 wbs_ufp_adr_i[6]
port 177 nsew signal input
rlabel metal3 s 11200 12248 12000 12368 6 wbs_ufp_adr_i[7]
port 178 nsew signal input
rlabel metal3 s 11200 13064 12000 13184 6 wbs_ufp_adr_i[8]
port 179 nsew signal input
rlabel metal3 s 11200 13744 12000 13864 6 wbs_ufp_adr_i[9]
port 180 nsew signal input
rlabel metal3 s 11200 2456 12000 2576 6 wbs_ufp_cyc_i
port 181 nsew signal input
rlabel metal3 s 11200 31152 12000 31272 6 wbs_ufp_dat_i[0]
port 182 nsew signal input
rlabel metal3 s 11200 38632 12000 38752 6 wbs_ufp_dat_i[10]
port 183 nsew signal input
rlabel metal3 s 11200 39448 12000 39568 6 wbs_ufp_dat_i[11]
port 184 nsew signal input
rlabel metal3 s 11200 40264 12000 40384 6 wbs_ufp_dat_i[12]
port 185 nsew signal input
rlabel metal3 s 11200 40944 12000 41064 6 wbs_ufp_dat_i[13]
port 186 nsew signal input
rlabel metal3 s 11200 41760 12000 41880 6 wbs_ufp_dat_i[14]
port 187 nsew signal input
rlabel metal3 s 11200 42440 12000 42560 6 wbs_ufp_dat_i[15]
port 188 nsew signal input
rlabel metal3 s 11200 43256 12000 43376 6 wbs_ufp_dat_i[16]
port 189 nsew signal input
rlabel metal3 s 11200 43936 12000 44056 6 wbs_ufp_dat_i[17]
port 190 nsew signal input
rlabel metal3 s 11200 44752 12000 44872 6 wbs_ufp_dat_i[18]
port 191 nsew signal input
rlabel metal3 s 11200 45432 12000 45552 6 wbs_ufp_dat_i[19]
port 192 nsew signal input
rlabel metal3 s 11200 31832 12000 31952 6 wbs_ufp_dat_i[1]
port 193 nsew signal input
rlabel metal3 s 11200 46248 12000 46368 6 wbs_ufp_dat_i[20]
port 194 nsew signal input
rlabel metal3 s 11200 46928 12000 47048 6 wbs_ufp_dat_i[21]
port 195 nsew signal input
rlabel metal3 s 11200 47744 12000 47864 6 wbs_ufp_dat_i[22]
port 196 nsew signal input
rlabel metal3 s 11200 48560 12000 48680 6 wbs_ufp_dat_i[23]
port 197 nsew signal input
rlabel metal3 s 11200 49240 12000 49360 6 wbs_ufp_dat_i[24]
port 198 nsew signal input
rlabel metal3 s 11200 50056 12000 50176 6 wbs_ufp_dat_i[25]
port 199 nsew signal input
rlabel metal3 s 11200 50736 12000 50856 6 wbs_ufp_dat_i[26]
port 200 nsew signal input
rlabel metal3 s 11200 51552 12000 51672 6 wbs_ufp_dat_i[27]
port 201 nsew signal input
rlabel metal3 s 11200 52232 12000 52352 6 wbs_ufp_dat_i[28]
port 202 nsew signal input
rlabel metal3 s 11200 53048 12000 53168 6 wbs_ufp_dat_i[29]
port 203 nsew signal input
rlabel metal3 s 11200 32648 12000 32768 6 wbs_ufp_dat_i[2]
port 204 nsew signal input
rlabel metal3 s 11200 53728 12000 53848 6 wbs_ufp_dat_i[30]
port 205 nsew signal input
rlabel metal3 s 11200 54544 12000 54664 6 wbs_ufp_dat_i[31]
port 206 nsew signal input
rlabel metal3 s 11200 33464 12000 33584 6 wbs_ufp_dat_i[3]
port 207 nsew signal input
rlabel metal3 s 11200 34144 12000 34264 6 wbs_ufp_dat_i[4]
port 208 nsew signal input
rlabel metal3 s 11200 34960 12000 35080 6 wbs_ufp_dat_i[5]
port 209 nsew signal input
rlabel metal3 s 11200 35640 12000 35760 6 wbs_ufp_dat_i[6]
port 210 nsew signal input
rlabel metal3 s 11200 36456 12000 36576 6 wbs_ufp_dat_i[7]
port 211 nsew signal input
rlabel metal3 s 11200 37136 12000 37256 6 wbs_ufp_dat_i[8]
port 212 nsew signal input
rlabel metal3 s 11200 37952 12000 38072 6 wbs_ufp_dat_i[9]
port 213 nsew signal input
rlabel metal3 s 11200 56040 12000 56160 6 wbs_ufp_dat_o[0]
port 214 nsew signal tristate
rlabel metal3 s 11200 63520 12000 63640 6 wbs_ufp_dat_o[10]
port 215 nsew signal tristate
rlabel metal3 s 11200 64336 12000 64456 6 wbs_ufp_dat_o[11]
port 216 nsew signal tristate
rlabel metal3 s 11200 65152 12000 65272 6 wbs_ufp_dat_o[12]
port 217 nsew signal tristate
rlabel metal3 s 11200 65832 12000 65952 6 wbs_ufp_dat_o[13]
port 218 nsew signal tristate
rlabel metal3 s 11200 66648 12000 66768 6 wbs_ufp_dat_o[14]
port 219 nsew signal tristate
rlabel metal3 s 11200 67328 12000 67448 6 wbs_ufp_dat_o[15]
port 220 nsew signal tristate
rlabel metal3 s 11200 68144 12000 68264 6 wbs_ufp_dat_o[16]
port 221 nsew signal tristate
rlabel metal3 s 11200 68824 12000 68944 6 wbs_ufp_dat_o[17]
port 222 nsew signal tristate
rlabel metal3 s 11200 69640 12000 69760 6 wbs_ufp_dat_o[18]
port 223 nsew signal tristate
rlabel metal3 s 11200 70320 12000 70440 6 wbs_ufp_dat_o[19]
port 224 nsew signal tristate
rlabel metal3 s 11200 56856 12000 56976 6 wbs_ufp_dat_o[1]
port 225 nsew signal tristate
rlabel metal3 s 11200 71136 12000 71256 6 wbs_ufp_dat_o[20]
port 226 nsew signal tristate
rlabel metal3 s 11200 71816 12000 71936 6 wbs_ufp_dat_o[21]
port 227 nsew signal tristate
rlabel metal3 s 11200 72632 12000 72752 6 wbs_ufp_dat_o[22]
port 228 nsew signal tristate
rlabel metal3 s 11200 73448 12000 73568 6 wbs_ufp_dat_o[23]
port 229 nsew signal tristate
rlabel metal3 s 11200 74128 12000 74248 6 wbs_ufp_dat_o[24]
port 230 nsew signal tristate
rlabel metal3 s 11200 74944 12000 75064 6 wbs_ufp_dat_o[25]
port 231 nsew signal tristate
rlabel metal3 s 11200 75624 12000 75744 6 wbs_ufp_dat_o[26]
port 232 nsew signal tristate
rlabel metal3 s 11200 76440 12000 76560 6 wbs_ufp_dat_o[27]
port 233 nsew signal tristate
rlabel metal3 s 11200 77120 12000 77240 6 wbs_ufp_dat_o[28]
port 234 nsew signal tristate
rlabel metal3 s 11200 77936 12000 78056 6 wbs_ufp_dat_o[29]
port 235 nsew signal tristate
rlabel metal3 s 11200 57536 12000 57656 6 wbs_ufp_dat_o[2]
port 236 nsew signal tristate
rlabel metal3 s 11200 78616 12000 78736 6 wbs_ufp_dat_o[30]
port 237 nsew signal tristate
rlabel metal3 s 11200 79432 12000 79552 6 wbs_ufp_dat_o[31]
port 238 nsew signal tristate
rlabel metal3 s 11200 58352 12000 58472 6 wbs_ufp_dat_o[3]
port 239 nsew signal tristate
rlabel metal3 s 11200 59032 12000 59152 6 wbs_ufp_dat_o[4]
port 240 nsew signal tristate
rlabel metal3 s 11200 59848 12000 59968 6 wbs_ufp_dat_o[5]
port 241 nsew signal tristate
rlabel metal3 s 11200 60528 12000 60648 6 wbs_ufp_dat_o[6]
port 242 nsew signal tristate
rlabel metal3 s 11200 61344 12000 61464 6 wbs_ufp_dat_o[7]
port 243 nsew signal tristate
rlabel metal3 s 11200 62024 12000 62144 6 wbs_ufp_dat_o[8]
port 244 nsew signal tristate
rlabel metal3 s 11200 62840 12000 62960 6 wbs_ufp_dat_o[9]
port 245 nsew signal tristate
rlabel metal3 s 11200 3952 12000 4072 6 wbs_ufp_sel_i[0]
port 246 nsew signal input
rlabel metal3 s 11200 4768 12000 4888 6 wbs_ufp_sel_i[1]
port 247 nsew signal input
rlabel metal3 s 11200 5448 12000 5568 6 wbs_ufp_sel_i[2]
port 248 nsew signal input
rlabel metal3 s 11200 6264 12000 6384 6 wbs_ufp_sel_i[3]
port 249 nsew signal input
rlabel metal3 s 11200 1776 12000 1896 6 wbs_ufp_stb_i
port 250 nsew signal input
rlabel metal3 s 11200 3272 12000 3392 6 wbs_ufp_we_i
port 251 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12000 80000
<< end >>
